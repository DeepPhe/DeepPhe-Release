Default Paragraph||(?:(?:[\t ]*\r?\n){2,})
Numbered Part||(?:\r?\n(?=PARTS?\s+\d+(?:\s+AND\s+\d+)?:))$
Section Part||(?:^[\t ]*PART[\t ]+\d+[^\n]*\n)
