-geographically determined (yes/no)|*patient ID|cancer link|*body location|body location laterality|body location clockface position|body location quadrant|Diagnosis|tumor type|cancer type|histologic type|tumor extent|er status interpretation|er status numeric value|er status method|pr status interpretation|pr status numeric value|pr status method|her2neu status interpretation|her2neu status numeric value|her2neu status method|radiologic tumor size (mm)|radiologic tumor size procedure method|pathologic tumor size (mm)|pathologic aggregate tumor size (mm)|calcificationsYes|patientX|cancer_patientX_Left_Breast_Current|Breast|Left|10_30_o_clock_position|Upper_Outer_Quadrant_of_the_Breast|Invasive_Ductal_Carcinoma_Not_Otherwise_Specified|PrimaryTumor|Adenocarcinoma|Ductal|Invasive_Lesion|Negative|0|Immunohistochemical_Test|Negative|0|Immunohistochemical_Test|Negative|0|Immunohistochemical_Test|12X34X56|Ultrasonography|13||PresentYes|patientX|cancer_patientX_Left_Breast_Current|Axillary_Lymph_Node|Left|||Metastatic_Carcinoma|Regional_Metastasis|Adenocarcinoma||||||||||||||||Absent