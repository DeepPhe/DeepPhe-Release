// TODO  - Rewrite with ontology sites.
// Add A "Major" site since .0 isn't always what we want.
//    e.g. Colon, NOS is C18.9 - while C18.0 is Appendix, which is not the major site.
// Use an asterisk   C18*|Colon

C000|Lip_Proper
C001|Lip_Proper
C002|Lip_Proper
C003|Lip_Proper
C004|Lip_Proper
C005|Lip_Proper
C006|Lip_Proper
C008|Lip_Proper
C009|Lip_Proper

C019|Root_Of_Tongue
C02*|Tongue
C020|Dorsal_Surface_Of_Tongue
C021|Border_Of_Tongue
C022|Ventral_Surface_Of_Tongue_NOS
C023|Body_Of_Tongue
C024|Lingual_Tonsil
C028|Junctional_Zone_Of_Tongue
C029|Tongue

C030|Sublingual_Region
C031|Sublingual_Region
C039|Sublingual_Region
C040|Sublingual_Region
C041|Sublingual_Region
C048|Sublingual_Region
C049|Sublingual_Region
C050|Sublingual_Region
C051|Sublingual_Region
C052|Sublingual_Region
C058|Sublingual_Region
C059|Sublingual_Region
C060|Sublingual_Region
C061|Sublingual_Region
C062|Sublingual_Region
C068|Sublingual_Region
C069|Sublingual_Region

C079|Salivary_Gland
C080|Salivary_Gland
C081|Salivary_Gland
C088|Salivary_Gland
C089|Salivary_Gland

// Actually Oropharynx.  Pharynx is C14*
C090|Pharynx
C091|Pharynx
C098|Pharynx
C099|Pharynx
C100|Pharynx
C101|Pharynx
C102|Pharynx
C103|Pharynx
C104|Pharynx
C108|Pharynx
C109|Pharynx

C110|Nasopharynx
C112|Nasopharynx
C113|Nasopharynx
C118|Nasopharynx
C119|Nasopharynx
C111|Posterior_Wall_Of_The_Nasopharynx

C129|Hypopharynx
C130|Hypopharynx
C131|Hypopharynx
C132|Hypopharynx
C138|Hypopharynx
C139|Hypopharynx

C140|Pharynx
C142|Pharynx
C148|Pharynx

C150|Esophagus
C151|Esophagus
C152|Esophagus
C153|Esophagus
C154|Esophagus
C155|Esophagus
C158|Esophagus
C159|Esophagus

C160|Stomach
C161|Stomach
C162|Stomach
C163|Stomach
C164|Stomach
C165|Stomach
C166|Stomach
C168|Stomach
C169|Stomach

C170|Duodenum
C171|Jejunum
C172|Ileum
C173|Meckel_Diverticulum
C178|Overlapping_Lesion_Of_Small_Intestine
C179|Small_Intestine

C18*|Colon
C180|Cecum
C181|Appendix
C182|Ascending_Colon
C183|Hepatic_Flexure
C184|Transverse_Colon
C185|Splenic_Flexure
// C186 in ontology is Left_Colon aka Descending_Colon
C186|Large_Intestine
C187|Sigmoid_Colon
C188|Overlapping_Lesion_Of_Colon
C189|Large_Intestine

C190|Rectosigmoid_Colon
C199|Rectosigmoid_Colon

C200|Rectal
C209|Rectal

C210|Anus
C211|Anal_Sphincter
C212|Cloacogenic_Zone
C218|Anorectal_Junction

C220|Liver
C221|Intrahepatic_Bile_Duct

// Actually Gall Bladder and Extrahepatic Bile Ducts
C239|Extrahepatic_Bile_Duct

C240|Extrahepatic_Bile_Duct
C241|Extrahepatic_Bile_Duct
C248|Extrahepatic_Bile_Duct
C249|Extrahepatic_Bile_Duct

C250|Pancreas
C251|Pancreas
C252|Pancreas
C253|Pancreas
C254|Pancreas
C257|Pancreas
C258|Pancreas
C259|Pancreas

// Actually Unspecified Digestive Organ
C260|Intestine
// C268 in ontology is (old) Overlapping_Lesion_Of_Digestive_System
C268|Overlapping_Lesion_Of_Digestive_System
// C269 in ontology is Entire_Digestive_Organ and ancestor Gastrointestinal_System
C269|Entire_Digestive_Organ
// Actually Nasal Cavity (including Nasal Cartilage)
// In Ontology is Nasal_Cavity and subclasses, including Nasal_Cartilage

C300|Nasal_Cartilage
C301|Middle_Ear

C310|Nasal_Sinus
C311|Nasal_Sinus
C312|Nasal_Sinus
C313|Nasal_Sinus
C318|Nasal_Sinus
// Actually Accessory Sinus, NOS
C319|Nasal_Sinus

C320|Larynx
C321|Larynx
C322|Larynx
C323|Larynx
C328|Larynx
C329|Larynx

C339|Trachea

// Actually Lung and Bronchus
C340|Bronchus
C341|Bronchus
C342|Bronchus
C343|Bronchus
C348|Bronchus
C349|Bronchus

C379|Thymus_Gland

C380|Heart
C381|Mediastinum
C382|Mediastinum
C383|Mediastinum
C384|Pleura
C388|Mediastinum

C390|Respiratory_System
C398|Respiratory_System
C399|Respiratory_System

// Should be Bones & Joints, excluding Skull, bones of face and mandible!
C400|Mandible
C401|Mandible
C402|Mandible
C403|Mandible
C408|Mandible
C409|Mandible

C410|Skull
C411|Mandible
C412|Mandible
C413|Mandible
C414|Mandible
C418|Mandible
C419|Mandible

// Actually Blood, Bone Marrow and Hematopoietic system
C420|Bone_Marrow
C421|Bone_Marrow
C422|Spleen
C423|Reticuloendothelial_System
C424|Bone_Marrow

C440|Skin
C441|Skin
C442|Skin
C443|Skin
C444|Skin
C445|Skin
C446|Skin
C447|Skin
C448|Skin
C449|Skin

C470|Peripheral_Nerve
C471|Peripheral_Nerve
C472|Peripheral_Nerve
C473|Peripheral_Nerve
C474|Peripheral_Nerve
C475|Peripheral_Nerve
C476|Peripheral_Nerve
C478|Peripheral_Nerve
C479|Peripheral_Nerve

// Actually Retroperitoneum and Peritoneum
C480|Retroperitoneal_Space
C481|Retroperitoneal_Space
C482|Retroperitoneal_Space
C488|Retroperitoneal_Space

// Actually Connective and Soft Tissue
C490|Body_Tissue
C491|Body_Tissue
C492|Body_Tissue
C493|Body_Tissue
C494|Body_Tissue
C495|Body_Tissue
C496|Body_Tissue
C498|Body_Tissue
C499|Body_Tissue

C50*|Breast
//C500|Nipple
C500|Breast
C501|Breast
C502|Upper_Inner_Quadrant
C503|Lower_Inner_Quadrant
C504|Upper_Outer_Quadrant
C505|Lower_Outer_Quadrant
C506|Breast
C508|Breast
C509|Breast

// Actually Vagina and Labia
C510|Vagina
C511|Vagina
C512|Vagina
C518|Vagina
C519|Vulva

C520|Vagina
C529|Vagina

C530|Cervix_Uteri
C531|Cervix_Uteri
C538|Cervix_Uteri
C539|Cervix_Uteri
C540|Corpus_Uteri
C541|Corpus_Uteri
C542|Corpus_Uteri
C543|Corpus_Uteri
C548|Corpus_Uteri
C549|Corpus_Uteri

C559|Uterus

C560|Ovary
C569|Ovary

C570|Fallopian_Tube
// Should be Other Female Genitalia excluding Fallopian Tube
C571|Fallopian_Tube
C572|Fallopian_Tube
C573|Fallopian_Tube
C574|Fallopian_Tube
C577|Fallopian_Tube
C578|Fallopian_Tube
C579|Fallopian_Tube

C589|Placenta_Part

C600|Penis
C601|Penis
C602|Penis
C608|Penis
C609|Penis

C610|Prostate
C619|Prostate

C620|Testis
C621|Testis
C629|Testis

// Actually Epididymis, Sperm Cord and Male Genitals NOS
C630|Spermatic_Cord
C631|Spermatic_Cord
C632|Scrotum
C637|Spermatic_Cord
C638|Spermatic_Cord
C639|Spermatic_Cord

C640|Kidney
C649|Kidney

// Actually Renal Pelvis, Ureter
C650|Pelvis
C659|Renal_Pelvis

C660|Pelvis
C669|Renal_Pelvis

C670|Urinary_Bladder
C671|Urinary_Bladder
C672|Urinary_Bladder
C673|Urinary_Bladder
C674|Urinary_Bladder
C675|Urinary_Bladder
C676|Urinary_Bladder
C677|Urinary_Bladder
C678|Urinary_Bladder
C679|Urinary_Bladder

// Actually Other Urinary Organs
C680|Genitourinary_System
C681|Genitourinary_System
C688|Genitourinary_System
C689|Genitourinary_System

// Actually Orbit and Lacrimal Gland
C690|Lacrimal_Gland
C691|Lacrimal_Gland
C692|Retina
C693|Lacrimal_Gland
// Actually Eyeball
C694|Eye
C695|Lacrimal_Gland
C696|Lacrimal_Gland
C697|Lacrimal_Gland
C698|Lacrimal_Gland
// Actually Eye, NOS
C699|Eye

C700|Meninges
C701|Meninges
C709|Meninges

// Should be Brain, Cranial Nerves and Spinal Cord
C710|Cranial_Nerve
C711|Cranial_Nerve
C712|Cranial_Nerve
C713|Cranial_Nerve
C714|Cranial_Nerve
C715|Heart_Ventricle
C716|Cerebellum
C717|Cranial_Nerve
C718|Cranial_Nerve
C719|Cranial_Nerve

C720|Cranial_Nerve
C721|Cranial_Nerve
C722|Cranial_Nerve
C723|Cranial_Nerve
C724|Cranial_Nerve
C725|Cranial_Nerve
// Other Nervous System
C728|Central_Nervous_System
C729|Central_Nervous_System

C730|Thyroid_Gland
C739|Thyroid_Gland

C740|Adrenal_Gland
C741|Adrenal_Gland
C749|Adrenal_Gland

C750|Parathyroid_Gland
C751|Pituitary_Gland
C752|Craniopharyngeal_Duct
C753|Pineal_Gland
// Actually Other Endocrine Glands
C754|Endocrine_Gland
C755|Endocrine_Gland
C758|Endocrine_Gland
C759|Endocrine_Gland

// Actually "Ill-Defined"
C760|Body_Region
C761|Body_Region
C762|Body_Region
C763|Body_Region
C764|Body_Region
C765|Body_Region
C766|Body_Region
C767|Body_Region
C768|Body_Region

C770|Lymph_Node
C771|Lymph_Node
C772|Lymph_Node
C773|Lymph_Node
C774|Lymph_Node
C775|Lymph_Node
C778|Lymph_Node
C779|Lymph_Node

C809|Undetermined
