Blank Line||(?:(?:\r?\n){2,})
Numbered Part||(?:\r?\n(?=PARTS?\s+\d+(?:\s+AND\s+\d+)?:))
