Default Paragraph||^[\t ]*\r?\n
//Numbered Part||(?:\r?\n(?=PARTS?\s+\d+(?:\s+AND\s+\d+)?:))$
//Section Part||(?:^[\t ]*PART[\t ]+\d+[^\n]*\n)
Dash Separator||^[\t ]*[-_=]{3,}[\t ]*\r?\n||^[\t ]*[-_=]{3,}[\t ]*\r?\n
