C800|Undetermined|850|DuctalCarcinoma|8500/1|DuctalCarcinoma
C800|Undetermined|807|SquamousCellNeoplasm|8070/1|SquamousCellNeoplasm
C000-C006,C008-C009|LipProper|801|Carcinoma|8010/2|InSituCancer
C000-C006,C008-C009|LipProper|801|Carcinoma|8010/3|CarcinomaNOSDNE
C000-C006,C008-C009|LipProper|801|Carcinoma|8011/3|MalignantEpithelioma
C000-C006,C008-C009|LipProper|801|Carcinoma|8012/3|LargeCellCarcinoma
C000-C006,C008-C009|LipProper|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C000-C006,C008-C009|LipProper|801|Carcinoma|8014/3|LargeCellCarcinoma
C000-C006,C008-C009|LipProper|801|Carcinoma|8015/3|GlassyCellCarcinoma
C000-C006,C008-C009|LipProper|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C000-C006,C008-C009|LipProper|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C000-C006,C008-C009|LipProper|802|Carcinoma|8022/3|PleomorphicCarcinoma
C000-C006,C008-C009|LipProper|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C000-C006,C008-C009|LipProper|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C000-C006,C008-C009|LipProper|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C000-C006,C008-C009|LipProper|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C000-C006,C008-C009|LipProper|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C000-C006,C008-C009|LipProper|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C000-C006,C008-C009|LipProper|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C000-C006,C008-C009|LipProper|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C000-C006,C008-C009|LipProper|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C000-C006,C008-C009|LipProper|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C000-C006,C008-C009|LipProper|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C000-C006,C008-C009|LipProper|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C000-C006,C008-C009|LipProper|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C000-C006,C008-C009|LipProper|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C000-C006,C008-C009|LipProper|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C000-C006,C008-C009|LipProper|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C000-C006,C008-C009|LipProper|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C000-C006,C008-C009|LipProper|814|Adenocarcinoma|8140/3|Adenocarcinoma
C000-C006,C008-C009|LipProper|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C000-C006,C008-C009|LipProper|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C000-C006,C008-C009|LipProper|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C000-C006,C008-C009|LipProper|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C000-C006,C008-C009|LipProper|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C000-C006,C008-C009|LipProper|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C000-C006,C008-C009|LipProper|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C000-C006,C008-C009|LipProper|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C000-C006,C008-C009|LipProper|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C000-C006,C008-C009|LipProper|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C000-C006,C008-C009|LipProper|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C000-C006,C008-C009|LipProper|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C000-C006,C008-C009|LipProper|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C000-C006,C008-C009|LipProper|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C000-C006,C008-C009|LipProper|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C000-C006,C008-C009|LipProper|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C000-C006,C008-C009|LipProper|872|Melanoma|8720/2|Stage0SkinMelanoma
C000-C006,C008-C009|LipProper|872|Melanoma|8720/3|Melanoma
C000-C006,C008-C009|LipProper|872|Melanoma|8721/3|NodularMelanoma
C000-C006,C008-C009|LipProper|872|Melanoma|8722/3|BalloonCellMelanoma
C000-C006,C008-C009|LipProper|872|Melanoma|8723/3|RegressingMelanoma
C000-C006,C008-C009|LipProper|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C000-C006,C008-C009|LipProper|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C000-C006,C008-C009|LipProper|874|Nevus|8745/3|DesmoplasticMelanoma
C000-C006,C008-C009|LipProper|874|Nevus|8746/3|MucosalLentiginousMelanoma
C000-C006,C008-C009|LipProper|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C000-C006,C008-C009|LipProper|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C000-C006,C008-C009|LipProper|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C000-C006,C008-C009|LipProper|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C000-C006,C008-C009|LipProper|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C000-C006,C008-C009|LipProper|914|KaposiSarcoma|9140/3|KaposiSarcoma
C000-C006,C008-C009|LipProper|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C000-C006,C008-C009|LipProper|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C019|RootOfTongue|801|Carcinoma|8010/2|InSituCancer
C019|RootOfTongue|801|Carcinoma|8010/3|CarcinomaNOSDNE
C019|RootOfTongue|801|Carcinoma|8011/3|MalignantEpithelioma
C019|RootOfTongue|801|Carcinoma|8012/3|LargeCellCarcinoma
C019|RootOfTongue|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C019|RootOfTongue|801|Carcinoma|8014/3|LargeCellCarcinoma
C019|RootOfTongue|801|Carcinoma|8015/3|GlassyCellCarcinoma
C019|RootOfTongue|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C019|RootOfTongue|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C019|RootOfTongue|802|Carcinoma|8022/3|PleomorphicCarcinoma
C019|RootOfTongue|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C019|RootOfTongue|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C019|RootOfTongue|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C019|RootOfTongue|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C019|RootOfTongue|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C019|RootOfTongue|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C019|RootOfTongue|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C019|RootOfTongue|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C019|RootOfTongue|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C019|RootOfTongue|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C019|RootOfTongue|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C019|RootOfTongue|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C019|RootOfTongue|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C019|RootOfTongue|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C019|RootOfTongue|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C019|RootOfTongue|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C019|RootOfTongue|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C019|RootOfTongue|808|LymphoepithelialCarcinoma|8085/3|SquamousCellCarcinoma
C019|RootOfTongue|808|LymphoepithelialCarcinoma|8086/3|SquamousCellCarcinoma
C019|RootOfTongue|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C019|RootOfTongue|814|Adenocarcinoma|8140/3|Adenocarcinoma
C019|RootOfTongue|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C019|RootOfTongue|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C019|RootOfTongue|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C019|RootOfTongue|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C019|RootOfTongue|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C019|RootOfTongue|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C019|RootOfTongue|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C019|RootOfTongue|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C019|RootOfTongue|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C019|RootOfTongue|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C019|RootOfTongue|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C019|RootOfTongue|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C019|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C019|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C019|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCellSpindleCell
C019|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C019|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C019|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C019|RootOfTongue|872|Melanoma|8720/2|Stage0SkinMelanoma
C019|RootOfTongue|872|Melanoma|8720/3|Melanoma
C019|RootOfTongue|872|Melanoma|8721/3|NodularMelanoma
C019|RootOfTongue|872|Melanoma|8722/3|BalloonCellMelanoma
C019|RootOfTongue|872|Melanoma|8723/3|RegressingMelanoma
C019|RootOfTongue|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C019|RootOfTongue|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C019|RootOfTongue|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C019|RootOfTongue|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C019|RootOfTongue|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C019|RootOfTongue|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C019|RootOfTongue|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C019|RootOfTongue|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C019|RootOfTongue|914|KaposiSarcoma|9140/3|KaposiSarcoma
C019|RootOfTongue|959|Lymphoma|9590/3|Lymphoma
C019|RootOfTongue|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C019|RootOfTongue|959|Lymphoma|9596/3|CompositeLymphoma
C019|RootOfTongue|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C019|RootOfTongue|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C019|RootOfTongue|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C019|RootOfTongue|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C019|RootOfTongue|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C019|RootOfTongue|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C019|RootOfTongue|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C019|RootOfTongue|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C019|RootOfTongue|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C019|RootOfTongue|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C019|RootOfTongue|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C019|RootOfTongue|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C019|RootOfTongue|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C019|RootOfTongue|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C019|RootOfTongue|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C019|RootOfTongue|967|BCellLymphomas|9673/3|MantleCellLymphoma
C019|RootOfTongue|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C019|RootOfTongue|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C019|RootOfTongue|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C019|RootOfTongue|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C019|RootOfTongue|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C019|RootOfTongue|969|FollicularAdenoma|9690/3|LymphomaFollicular
C019|RootOfTongue|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C019|RootOfTongue|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C019|RootOfTongue|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C019|RootOfTongue|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C019|RootOfTongue|970|TCellLymphoma|9701/3|SezarySyndrome
C019|RootOfTongue|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C019|RootOfTongue|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C019|RootOfTongue|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C019|RootOfTongue|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C019|RootOfTongue|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C019|RootOfTongue|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C019|RootOfTongue|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C019|RootOfTongue|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C019|RootOfTongue|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C019|RootOfTongue|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C019|RootOfTongue|973|Plasmacytoma|9731/3|Plasmacytoma
C019|RootOfTongue|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C019|RootOfTongue|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C019|RootOfTongue|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C019|RootOfTongue|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C019|RootOfTongue|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C019|RootOfTongue|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C019|RootOfTongue|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C019|RootOfTongue|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C019|RootOfTongue|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C019|RootOfTongue|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C019|RootOfTongue|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C019|RootOfTongue|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C019|RootOfTongue|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C019|RootOfTongue|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C019|RootOfTongue|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C019|RootOfTongue|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9812/3|null
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9813/3|null
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9814/3|null
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9817/3|null
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9818/3|null
C019|RootOfTongue|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C019|RootOfTongue|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C019|RootOfTongue|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C019|RootOfTongue|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C019|RootOfTongue|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C019|RootOfTongue|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C019|RootOfTongue|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C019|RootOfTongue|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C020-C024,C028-C029|RootOfTongue|801|Carcinoma|8010/2|InSituCancer
C020-C024,C028-C029|RootOfTongue|801|Carcinoma|8010/3|CarcinomaNOSDNE
C020-C024,C028-C029|RootOfTongue|801|Carcinoma|8011/3|MalignantEpithelioma
C020-C024,C028-C029|RootOfTongue|801|Carcinoma|8012/3|LargeCellCarcinoma
C020-C024,C028-C029|RootOfTongue|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C020-C024,C028-C029|RootOfTongue|801|Carcinoma|8014/3|LargeCellCarcinoma
C020-C024,C028-C029|RootOfTongue|801|Carcinoma|8015/3|GlassyCellCarcinoma
C020-C024,C028-C029|RootOfTongue|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C020-C024,C028-C029|RootOfTongue|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C020-C024,C028-C029|RootOfTongue|802|Carcinoma|8022/3|PleomorphicCarcinoma
C020-C024,C028-C029|RootOfTongue|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C020-C024,C028-C029|RootOfTongue|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C020-C024,C028-C029|RootOfTongue|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C020-C024,C028-C029|RootOfTongue|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C020-C024,C028-C029|RootOfTongue|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C020-C024,C028-C029|RootOfTongue|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C020-C024,C028-C029|RootOfTongue|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C020-C024,C028-C029|RootOfTongue|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C020-C024,C028-C029|RootOfTongue|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C020-C024,C028-C029|RootOfTongue|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C020-C024,C028-C029|RootOfTongue|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C020-C024,C028-C029|RootOfTongue|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C020-C024,C028-C029|RootOfTongue|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C020-C024,C028-C029|RootOfTongue|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C020-C024,C028-C029|RootOfTongue|814|Adenocarcinoma|8140/3|Adenocarcinoma
C020-C024,C028-C029|RootOfTongue|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C020-C024,C028-C029|RootOfTongue|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C020-C024,C028-C029|RootOfTongue|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C020-C024,C028-C029|RootOfTongue|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C020-C024,C028-C029|RootOfTongue|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C020-C024,C028-C029|RootOfTongue|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C020-C024,C028-C029|RootOfTongue|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C020-C024,C028-C029|RootOfTongue|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C020-C024,C028-C029|RootOfTongue|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C020-C024,C028-C029|RootOfTongue|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C020-C024,C028-C029|RootOfTongue|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C020-C024,C028-C029|RootOfTongue|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C020-C024,C028-C029|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C020-C024,C028-C029|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C020-C024,C028-C029|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCellSpindleCell
C020-C024,C028-C029|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C020-C024,C028-C029|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C020-C024,C028-C029|RootOfTongue|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C020-C024,C028-C029|RootOfTongue|872|Melanoma|8720/2|Stage0SkinMelanoma
C020-C024,C028-C029|RootOfTongue|872|Melanoma|8720/3|Melanoma
C020-C024,C028-C029|RootOfTongue|872|Melanoma|8721/3|NodularMelanoma
C020-C024,C028-C029|RootOfTongue|872|Melanoma|8722/3|BalloonCellMelanoma
C020-C024,C028-C029|RootOfTongue|872|Melanoma|8723/3|RegressingMelanoma
C020-C024,C028-C029|RootOfTongue|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C020-C024,C028-C029|RootOfTongue|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C020-C024,C028-C029|RootOfTongue|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C020-C024,C028-C029|RootOfTongue|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C020-C024,C028-C029|RootOfTongue|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C020-C024,C028-C029|RootOfTongue|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C020-C024,C028-C029|RootOfTongue|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C020-C024,C028-C029|RootOfTongue|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C020-C024,C028-C029|RootOfTongue|914|KaposiSarcoma|9140/3|KaposiSarcoma
C020-C024,C028-C029|RootOfTongue|959|Lymphoma|9590/3|Lymphoma
C020-C024,C028-C029|RootOfTongue|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C020-C024,C028-C029|RootOfTongue|959|Lymphoma|9596/3|CompositeLymphoma
C020-C024,C028-C029|RootOfTongue|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C020-C024,C028-C029|RootOfTongue|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C020-C024,C028-C029|RootOfTongue|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C020-C024,C028-C029|RootOfTongue|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C020-C024,C028-C029|RootOfTongue|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C020-C024,C028-C029|RootOfTongue|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C020-C024,C028-C029|RootOfTongue|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C020-C024,C028-C029|RootOfTongue|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C020-C024,C028-C029|RootOfTongue|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C020-C024,C028-C029|RootOfTongue|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C020-C024,C028-C029|RootOfTongue|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C020-C024,C028-C029|RootOfTongue|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C020-C024,C028-C029|RootOfTongue|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C020-C024,C028-C029|RootOfTongue|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C020-C024,C028-C029|RootOfTongue|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C020-C024,C028-C029|RootOfTongue|967|BCellLymphomas|9673/3|MantleCellLymphoma
C020-C024,C028-C029|RootOfTongue|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C020-C024,C028-C029|RootOfTongue|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C020-C024,C028-C029|RootOfTongue|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C020-C024,C028-C029|RootOfTongue|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C020-C024,C028-C029|RootOfTongue|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C020-C024,C028-C029|RootOfTongue|969|FollicularAdenoma|9690/3|LymphomaFollicular
C020-C024,C028-C029|RootOfTongue|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C020-C024,C028-C029|RootOfTongue|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C020-C024,C028-C029|RootOfTongue|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C020-C024,C028-C029|RootOfTongue|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C020-C024,C028-C029|RootOfTongue|970|TCellLymphoma|9701/3|SezarySyndrome
C020-C024,C028-C029|RootOfTongue|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C020-C024,C028-C029|RootOfTongue|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C020-C024,C028-C029|RootOfTongue|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C020-C024,C028-C029|RootOfTongue|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C020-C024,C028-C029|RootOfTongue|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C020-C024,C028-C029|RootOfTongue|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C020-C024,C028-C029|RootOfTongue|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C020-C024,C028-C029|RootOfTongue|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C020-C024,C028-C029|RootOfTongue|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C020-C024,C028-C029|RootOfTongue|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C020-C024,C028-C029|RootOfTongue|973|Plasmacytoma|9731/3|Plasmacytoma
C020-C024,C028-C029|RootOfTongue|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C020-C024,C028-C029|RootOfTongue|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C020-C024,C028-C029|RootOfTongue|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C020-C024,C028-C029|RootOfTongue|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C020-C024,C028-C029|RootOfTongue|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C020-C024,C028-C029|RootOfTongue|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C020-C024,C028-C029|RootOfTongue|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C020-C024,C028-C029|RootOfTongue|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C020-C024,C028-C029|RootOfTongue|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C020-C024,C028-C029|RootOfTongue|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C020-C024,C028-C029|RootOfTongue|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C020-C024,C028-C029|RootOfTongue|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C020-C024,C028-C029|RootOfTongue|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C020-C024,C028-C029|RootOfTongue|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C020-C024,C028-C029|RootOfTongue|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C020-C024,C028-C029|RootOfTongue|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9812/3|null
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9813/3|null
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9814/3|null
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9817/3|null
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9818/3|null
C020-C024,C028-C029|RootOfTongue|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C020-C024,C028-C029|RootOfTongue|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C020-C024,C028-C029|RootOfTongue|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C020-C024,C028-C029|RootOfTongue|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C020-C024,C028-C029|RootOfTongue|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C020-C024,C028-C029|RootOfTongue|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C020-C024,C028-C029|RootOfTongue|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C020-C024,C028-C029|RootOfTongue|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|801|Carcinoma|8010/2|InSituCancer
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|801|Carcinoma|8010/3|CarcinomaNOSDNE
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|801|Carcinoma|8011/3|MalignantEpithelioma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|801|Carcinoma|8012/3|LargeCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|801|Carcinoma|8014/3|LargeCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|801|Carcinoma|8015/3|GlassyCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|802|Carcinoma|8022/3|PleomorphicCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|814|Adenocarcinoma|8140/3|Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|872|Melanoma|8720/2|Stage0SkinMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|872|Melanoma|8720/3|Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|872|Melanoma|8721/3|NodularMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|872|Melanoma|8722/3|BalloonCellMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|872|Melanoma|8723/3|RegressingMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|874|Nevus|8745/3|DesmoplasticMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|874|Nevus|8746/3|MucosalLentiginousMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|898|Carcinosarcoma|8980/3|Carcinosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|914|KaposiSarcoma|9140/3|KaposiSarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|959|Lymphoma|9590/3|Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|959|Lymphoma|9596/3|CompositeLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|967|BCellLymphomas|9673/3|MantleCellLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|969|FollicularAdenoma|9690/3|LymphomaFollicular
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|970|TCellLymphoma|9701/3|SezarySyndrome
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|973|Plasmacytoma|9731/3|Plasmacytoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9812/3|null
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9813/3|null
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9814/3|null
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9817/3|null
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9818/3|null
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|SublingualRegion|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C079-C081,C088-C089|SalivaryGland|801|Carcinoma|8010/2|InSituCancer
C079-C081,C088-C089|SalivaryGland|801|Carcinoma|8010/3|CarcinomaNOSDNE
C079-C081,C088-C089|SalivaryGland|801|Carcinoma|8011/3|MalignantEpithelioma
C079-C081,C088-C089|SalivaryGland|801|Carcinoma|8012/3|LargeCellCarcinoma
C079-C081,C088-C089|SalivaryGland|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C079-C081,C088-C089|SalivaryGland|801|Carcinoma|8014/3|LargeCellCarcinoma
C079-C081,C088-C089|SalivaryGland|801|Carcinoma|8015/3|GlassyCellCarcinoma
C079-C081,C088-C089|SalivaryGland|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C079-C081,C088-C089|SalivaryGland|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C079-C081,C088-C089|SalivaryGland|802|Carcinoma|8022/3|PleomorphicCarcinoma
C079-C081,C088-C089|SalivaryGland|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C079-C081,C088-C089|SalivaryGland|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C079-C081,C088-C089|SalivaryGland|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C079-C081,C088-C089|SalivaryGland|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C079-C081,C088-C089|SalivaryGland|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C079-C081,C088-C089|SalivaryGland|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C079-C081,C088-C089|SalivaryGland|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C079-C081,C088-C089|SalivaryGland|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C079-C081,C088-C089|SalivaryGland|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C079-C081,C088-C089|SalivaryGland|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C079-C081,C088-C089|SalivaryGland|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C079-C081,C088-C089|SalivaryGland|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C079-C081,C088-C089|SalivaryGland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C079-C081,C088-C089|SalivaryGland|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C079-C081,C088-C089|SalivaryGland|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C079-C081,C088-C089|SalivaryGland|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C079-C081,C088-C089|SalivaryGland|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C079-C081,C088-C089|SalivaryGland|823|SolidCarcinoma|8230/2|InSituCancer
C079-C081,C088-C089|SalivaryGland|823|SolidCarcinoma|8230/3|SolidCarcinoma
C079-C081,C088-C089|SalivaryGland|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C079-C081,C088-C089|SalivaryGland|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C079-C081,C088-C089|SalivaryGland|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C079-C081,C088-C089|SalivaryGland|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C079-C081,C088-C089|SalivaryGland|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C079-C081,C088-C089|SalivaryGland|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C079-C081,C088-C089|SalivaryGland|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C079-C081,C088-C089|SalivaryGland|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C079-C081,C088-C089|SalivaryGland|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C079-C081,C088-C089|SalivaryGland|850|DuctalCarcinoma|8500/3|InvasiveBreastCarcinoma
C079-C081,C088-C089|SalivaryGland|850|DuctalCarcinoma|8502/3|SecretoryBreastCarcinoma
C079-C081,C088-C089|SalivaryGland|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C079-C081,C088-C089|SalivaryGland|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C079-C081,C088-C089|SalivaryGland|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C079-C081,C088-C089|SalivaryGland|856|AdenosquamousCarcinoma|8561/3|Adenolymphoma
C079-C081,C088-C089|SalivaryGland|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C079-C081,C088-C089|SalivaryGland|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C079-C081,C088-C089|SalivaryGland|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C079-C081,C088-C089|SalivaryGland|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCellSpindleCell
C079-C081,C088-C089|SalivaryGland|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C079-C081,C088-C089|SalivaryGland|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C079-C081,C088-C089|SalivaryGland|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C079-C081,C088-C089|SalivaryGland|880|Sarcoma|8800/3|Sarcoma
C079-C081,C088-C089|SalivaryGland|880|Sarcoma|8801/3|SpindleCellSarcoma
C079-C081,C088-C089|SalivaryGland|880|Sarcoma|8802/3|GiantCellSarcoma
C079-C081,C088-C089|SalivaryGland|880|Sarcoma|8803/3|SmallCellSarcoma
C079-C081,C088-C089|SalivaryGland|880|Sarcoma|8804/3|SarcomaEpithelioid
C079-C081,C088-C089|SalivaryGland|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C079-C081,C088-C089|SalivaryGland|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C079-C081,C088-C089|SalivaryGland|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C079-C081,C088-C089|SalivaryGland|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C079-C081,C088-C089|SalivaryGland|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C079-C081,C088-C089|SalivaryGland|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C079-C081,C088-C089|SalivaryGland|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C079-C081,C088-C089|SalivaryGland|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C079-C081,C088-C089|SalivaryGland|884|Myxosarcoma|8840/3|Myxosarcoma
C079-C081,C088-C089|SalivaryGland|885|Liposarcoma|8850/3|Liposarcoma
C079-C081,C088-C089|SalivaryGland|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C079-C081,C088-C089|SalivaryGland|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C079-C081,C088-C089|SalivaryGland|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C079-C081,C088-C089|SalivaryGland|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C079-C081,C088-C089|SalivaryGland|885|Liposarcoma|8855/3|Liposarcoma
C079-C081,C088-C089|SalivaryGland|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C079-C081,C088-C089|SalivaryGland|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C079-C081,C088-C089|SalivaryGland|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C079-C081,C088-C089|SalivaryGland|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C079-C081,C088-C089|SalivaryGland|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C079-C081,C088-C089|SalivaryGland|889|MyomatousNeoplasm|8895/3|Myosarcoma
C079-C081,C088-C089|SalivaryGland|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C079-C081,C088-C089|SalivaryGland|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C079-C081,C088-C089|SalivaryGland|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C079-C081,C088-C089|SalivaryGland|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C079-C081,C088-C089|SalivaryGland|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C079-C081,C088-C089|SalivaryGland|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C079-C081,C088-C089|SalivaryGland|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C079-C081,C088-C089|SalivaryGland|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C079-C081,C088-C089|SalivaryGland|898|Carcinosarcoma|8980/3|Carcinosarcoma
C079-C081,C088-C089|SalivaryGland|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C079-C081,C088-C089|SalivaryGland|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C079-C081,C088-C089|SalivaryGland|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C079-C081,C088-C089|SalivaryGland|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C079-C081,C088-C089|SalivaryGland|914|KaposiSarcoma|9140/3|KaposiSarcoma
C079-C081,C088-C089|SalivaryGland|959|Lymphoma|9590/3|Lymphoma
C079-C081,C088-C089|SalivaryGland|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C079-C081,C088-C089|SalivaryGland|959|Lymphoma|9596/3|CompositeLymphoma
C079-C081,C088-C089|SalivaryGland|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C079-C081,C088-C089|SalivaryGland|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C079-C081,C088-C089|SalivaryGland|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C079-C081,C088-C089|SalivaryGland|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C079-C081,C088-C089|SalivaryGland|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C079-C081,C088-C089|SalivaryGland|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C079-C081,C088-C089|SalivaryGland|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C079-C081,C088-C089|SalivaryGland|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C079-C081,C088-C089|SalivaryGland|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C079-C081,C088-C089|SalivaryGland|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C079-C081,C088-C089|SalivaryGland|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C079-C081,C088-C089|SalivaryGland|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C079-C081,C088-C089|SalivaryGland|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C079-C081,C088-C089|SalivaryGland|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C079-C081,C088-C089|SalivaryGland|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C079-C081,C088-C089|SalivaryGland|967|BCellLymphomas|9673/3|MantleCellLymphoma
C079-C081,C088-C089|SalivaryGland|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C079-C081,C088-C089|SalivaryGland|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C079-C081,C088-C089|SalivaryGland|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C079-C081,C088-C089|SalivaryGland|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C079-C081,C088-C089|SalivaryGland|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C079-C081,C088-C089|SalivaryGland|969|FollicularAdenoma|9690/3|LymphomaFollicular
C079-C081,C088-C089|SalivaryGland|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C079-C081,C088-C089|SalivaryGland|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C079-C081,C088-C089|SalivaryGland|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C079-C081,C088-C089|SalivaryGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C079-C081,C088-C089|SalivaryGland|970|TCellLymphoma|9701/3|SezarySyndrome
C079-C081,C088-C089|SalivaryGland|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C079-C081,C088-C089|SalivaryGland|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C079-C081,C088-C089|SalivaryGland|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C079-C081,C088-C089|SalivaryGland|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C079-C081,C088-C089|SalivaryGland|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C079-C081,C088-C089|SalivaryGland|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C079-C081,C088-C089|SalivaryGland|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C079-C081,C088-C089|SalivaryGland|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C079-C081,C088-C089|SalivaryGland|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C079-C081,C088-C089|SalivaryGland|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C079-C081,C088-C089|SalivaryGland|973|Plasmacytoma|9731/3|Plasmacytoma
C079-C081,C088-C089|SalivaryGland|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C079-C081,C088-C089|SalivaryGland|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C079-C081,C088-C089|SalivaryGland|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C079-C081,C088-C089|SalivaryGland|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C079-C081,C088-C089|SalivaryGland|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C079-C081,C088-C089|SalivaryGland|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C079-C081,C088-C089|SalivaryGland|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C079-C081,C088-C089|SalivaryGland|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C079-C081,C088-C089|SalivaryGland|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C079-C081,C088-C089|SalivaryGland|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C079-C081,C088-C089|SalivaryGland|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C079-C081,C088-C089|SalivaryGland|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C079-C081,C088-C089|SalivaryGland|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C079-C081,C088-C089|SalivaryGland|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C079-C081,C088-C089|SalivaryGland|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C079-C081,C088-C089|SalivaryGland|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9812/3|null
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9813/3|null
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9814/3|null
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9817/3|null
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9818/3|null
C079-C081,C088-C089|SalivaryGland|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C079-C081,C088-C089|SalivaryGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C079-C081,C088-C089|SalivaryGland|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C079-C081,C088-C089|SalivaryGland|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C079-C081,C088-C089|SalivaryGland|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C079-C081,C088-C089|SalivaryGland|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C079-C081,C088-C089|SalivaryGland|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C079-C081,C088-C089|SalivaryGland|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8010/2|InSituCancer
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8010/3|CarcinomaNOSDNE
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8011/3|MalignantEpithelioma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8012/3|LargeCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8014/3|LargeCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8015/3|GlassyCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C090-C091,C098-C104,C108-C109|Pharynx|802|Carcinoma|8022/3|PleomorphicCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C090-C091,C098-C104,C108-C109|Pharynx|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C090-C091,C098-C104,C108-C109|Pharynx|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C090-C091,C098-C104,C108-C109|Pharynx|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|LymphoepithelialCarcinoma|8085/3|SquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|LymphoepithelialCarcinoma|8086/3|SquamousCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C090-C091,C098-C104,C108-C109|Pharynx|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C090-C091,C098-C104,C108-C109|Pharynx|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C090-C091,C098-C104,C108-C109|Pharynx|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C090-C091,C098-C104,C108-C109|Pharynx|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C090-C091,C098-C104,C108-C109|Pharynx|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C090-C091,C098-C104,C108-C109|Pharynx|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C090-C091,C098-C104,C108-C109|Pharynx|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8720/2|Stage0SkinMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8720/3|Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8721/3|NodularMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8722/3|BalloonCellMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8723/3|RegressingMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C090-C091,C098-C104,C108-C109|Pharynx|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|874|Nevus|8745/3|DesmoplasticMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|874|Nevus|8746/3|MucosalLentiginousMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|876|Nevus|8761/3|GiantCongenitalNevus
C090-C091,C098-C104,C108-C109|Pharynx|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8800/3|Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8801/3|SpindleCellSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8802/3|GiantCellSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8803/3|SmallCellSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8804/3|SarcomaEpithelioid
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8850/3|Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8855/3|Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C090-C091,C098-C104,C108-C109|Pharynx|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C090-C091,C098-C104,C108-C109|Pharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C090-C091,C098-C104,C108-C109|Pharynx|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C090-C091,C098-C104,C108-C109|Pharynx|914|KaposiSarcoma|9140/3|KaposiSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|959|Lymphoma|9590/3|Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|959|Lymphoma|9596/3|CompositeLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C090-C091,C098-C104,C108-C109|Pharynx|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C090-C091,C098-C104,C108-C109|Pharynx|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C090-C091,C098-C104,C108-C109|Pharynx|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C090-C091,C098-C104,C108-C109|Pharynx|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C090-C091,C098-C104,C108-C109|Pharynx|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C090-C091,C098-C104,C108-C109|Pharynx|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C090-C091,C098-C104,C108-C109|Pharynx|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C090-C091,C098-C104,C108-C109|Pharynx|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C090-C091,C098-C104,C108-C109|Pharynx|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C090-C091,C098-C104,C108-C109|Pharynx|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|967|BCellLymphomas|9673/3|MantleCellLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|969|FollicularAdenoma|9690/3|LymphomaFollicular
C090-C091,C098-C104,C108-C109|Pharynx|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C090-C091,C098-C104,C108-C109|Pharynx|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C090-C091,C098-C104,C108-C109|Pharynx|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|970|TCellLymphoma|9701/3|SezarySyndrome
C090-C091,C098-C104,C108-C109|Pharynx|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C090-C091,C098-C104,C108-C109|Pharynx|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C090-C091,C098-C104,C108-C109|Pharynx|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C090-C091,C098-C104,C108-C109|Pharynx|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C090-C091,C098-C104,C108-C109|Pharynx|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C090-C091,C098-C104,C108-C109|Pharynx|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C090-C091,C098-C104,C108-C109|Pharynx|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C090-C091,C098-C104,C108-C109|Pharynx|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C090-C091,C098-C104,C108-C109|Pharynx|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C090-C091,C098-C104,C108-C109|Pharynx|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C090-C091,C098-C104,C108-C109|Pharynx|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C090-C091,C098-C104,C108-C109|Pharynx|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C090-C091,C098-C104,C108-C109|Pharynx|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9812/3|null
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9813/3|null
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9814/3|null
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9817/3|null
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9818/3|null
C090-C091,C098-C104,C108-C109|Pharynx|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C090-C091,C098-C104,C108-C109|Pharynx|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C090-C091,C098-C104,C108-C109|Pharynx|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C090-C091,C098-C104,C108-C109|Pharynx|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C090-C091,C098-C104,C108-C109|Pharynx|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C090-C091,C098-C104,C108-C109|Pharynx|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C090-C091,C098-C104,C108-C109|Pharynx|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C090-C091,C098-C104,C108-C109|Pharynx|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8010/2|InSituCancer
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8010/3|CarcinomaNOSDNE
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8011/3|MalignantEpithelioma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8012/3|LargeCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8014/3|LargeCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8015/3|GlassyCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C110,C112-C113,C118-C119|Nasopharynx|802|Carcinoma|8022/3|PleomorphicCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C110,C112-C113,C118-C119|Nasopharynx|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C110,C112-C113,C118-C119|Nasopharynx|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C110,C112-C113,C118-C119|Nasopharynx|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C110,C112-C113,C118-C119|Nasopharynx|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C110,C112-C113,C118-C119|Nasopharynx|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C110,C112-C113,C118-C119|Nasopharynx|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C110,C112-C113,C118-C119|Nasopharynx|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C110,C112-C113,C118-C119|Nasopharynx|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C110,C112-C113,C118-C119|Nasopharynx|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C110,C112-C113,C118-C119|Nasopharynx|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C110,C112-C113,C118-C119|Nasopharynx|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8720/2|Stage0SkinMelanoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8720/3|Melanoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8721/3|NodularMelanoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8722/3|BalloonCellMelanoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8723/3|RegressingMelanoma
C110,C112-C113,C118-C119|Nasopharynx|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C110,C112-C113,C118-C119|Nasopharynx|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C110,C112-C113,C118-C119|Nasopharynx|874|Nevus|8745/3|DesmoplasticMelanoma
C110,C112-C113,C118-C119|Nasopharynx|874|Nevus|8746/3|MucosalLentiginousMelanoma
C110,C112-C113,C118-C119|Nasopharynx|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C110,C112-C113,C118-C119|Nasopharynx|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C110,C112-C113,C118-C119|Nasopharynx|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8800/3|Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8801/3|SpindleCellSarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8802/3|GiantCellSarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8803/3|SmallCellSarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8804/3|SarcomaEpithelioid
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C110,C112-C113,C118-C119|Nasopharynx|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C110,C112-C113,C118-C119|Nasopharynx|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C110,C112-C113,C118-C119|Nasopharynx|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C110,C112-C113,C118-C119|Nasopharynx|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C110,C112-C113,C118-C119|Nasopharynx|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C110,C112-C113,C118-C119|Nasopharynx|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C110,C112-C113,C118-C119|Nasopharynx|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C110,C112-C113,C118-C119|Nasopharynx|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C110,C112-C113,C118-C119|Nasopharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C110,C112-C113,C118-C119|Nasopharynx|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C110,C112-C113,C118-C119|Nasopharynx|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C110,C112-C113,C118-C119|Nasopharynx|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C110,C112-C113,C118-C119|Nasopharynx|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C110,C112-C113,C118-C119|Nasopharynx|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C110,C112-C113,C118-C119|Nasopharynx|914|KaposiSarcoma|9140/3|KaposiSarcoma
C110,C112-C113,C118-C119|Nasopharynx|937|Chordoma|9370/3|Chordoma
C110,C112-C113,C118-C119|Nasopharynx|937|Chordoma|9371/3|ChondroidChordoma
C110,C112-C113,C118-C119|Nasopharynx|937|Chordoma|9372/3|DedifferentiatedChordoma
C110,C112-C113,C118-C119|Nasopharynx|959|Lymphoma|9590/3|Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C110,C112-C113,C118-C119|Nasopharynx|959|Lymphoma|9596/3|CompositeLymphoma
C110,C112-C113,C118-C119|Nasopharynx|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C110,C112-C113,C118-C119|Nasopharynx|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C110,C112-C113,C118-C119|Nasopharynx|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C110,C112-C113,C118-C119|Nasopharynx|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C110,C112-C113,C118-C119|Nasopharynx|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C110,C112-C113,C118-C119|Nasopharynx|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C110,C112-C113,C118-C119|Nasopharynx|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C110,C112-C113,C118-C119|Nasopharynx|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C110,C112-C113,C118-C119|Nasopharynx|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C110,C112-C113,C118-C119|Nasopharynx|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C110,C112-C113,C118-C119|Nasopharynx|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C110,C112-C113,C118-C119|Nasopharynx|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C110,C112-C113,C118-C119|Nasopharynx|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C110,C112-C113,C118-C119|Nasopharynx|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C110,C112-C113,C118-C119|Nasopharynx|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C110,C112-C113,C118-C119|Nasopharynx|967|BCellLymphomas|9673/3|MantleCellLymphoma
C110,C112-C113,C118-C119|Nasopharynx|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C110,C112-C113,C118-C119|Nasopharynx|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C110,C112-C113,C118-C119|Nasopharynx|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C110,C112-C113,C118-C119|Nasopharynx|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C110,C112-C113,C118-C119|Nasopharynx|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C110,C112-C113,C118-C119|Nasopharynx|969|FollicularAdenoma|9690/3|LymphomaFollicular
C110,C112-C113,C118-C119|Nasopharynx|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C110,C112-C113,C118-C119|Nasopharynx|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C110,C112-C113,C118-C119|Nasopharynx|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C110,C112-C113,C118-C119|Nasopharynx|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C110,C112-C113,C118-C119|Nasopharynx|970|TCellLymphoma|9701/3|SezarySyndrome
C110,C112-C113,C118-C119|Nasopharynx|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C110,C112-C113,C118-C119|Nasopharynx|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C110,C112-C113,C118-C119|Nasopharynx|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C110,C112-C113,C118-C119|Nasopharynx|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C110,C112-C113,C118-C119|Nasopharynx|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C110,C112-C113,C118-C119|Nasopharynx|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C110,C112-C113,C118-C119|Nasopharynx|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C110,C112-C113,C118-C119|Nasopharynx|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C110,C112-C113,C118-C119|Nasopharynx|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C110,C112-C113,C118-C119|Nasopharynx|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C110,C112-C113,C118-C119|Nasopharynx|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C110,C112-C113,C118-C119|Nasopharynx|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C110,C112-C113,C118-C119|Nasopharynx|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C110,C112-C113,C118-C119|Nasopharynx|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C110,C112-C113,C118-C119|Nasopharynx|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C110,C112-C113,C118-C119|Nasopharynx|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C110,C112-C113,C118-C119|Nasopharynx|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C110,C112-C113,C118-C119|Nasopharynx|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C110,C112-C113,C118-C119|Nasopharynx|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C110,C112-C113,C118-C119|Nasopharynx|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C110,C112-C113,C118-C119|Nasopharynx|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9812/3|null
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9813/3|null
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9814/3|null
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9817/3|null
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9818/3|null
C110,C112-C113,C118-C119|Nasopharynx|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C110,C112-C113,C118-C119|Nasopharynx|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C110,C112-C113,C118-C119|Nasopharynx|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C110,C112-C113,C118-C119|Nasopharynx|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C110,C112-C113,C118-C119|Nasopharynx|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C110,C112-C113,C118-C119|Nasopharynx|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C110,C112-C113,C118-C119|Nasopharynx|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C110,C112-C113,C118-C119|Nasopharynx|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C111|PosteriorWallOfTheNasopharynx|801|Carcinoma|8010/2|InSituCancer
C111|PosteriorWallOfTheNasopharynx|801|Carcinoma|8010/3|CarcinomaNOSDNE
C111|PosteriorWallOfTheNasopharynx|801|Carcinoma|8011/3|MalignantEpithelioma
C111|PosteriorWallOfTheNasopharynx|801|Carcinoma|8012/3|LargeCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C111|PosteriorWallOfTheNasopharynx|801|Carcinoma|8014/3|LargeCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|801|Carcinoma|8015/3|GlassyCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C111|PosteriorWallOfTheNasopharynx|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C111|PosteriorWallOfTheNasopharynx|802|Carcinoma|8022/3|PleomorphicCarcinoma
C111|PosteriorWallOfTheNasopharynx|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C111|PosteriorWallOfTheNasopharynx|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C111|PosteriorWallOfTheNasopharynx|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C111|PosteriorWallOfTheNasopharynx|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C111|PosteriorWallOfTheNasopharynx|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C111|PosteriorWallOfTheNasopharynx|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C111|PosteriorWallOfTheNasopharynx|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C111|PosteriorWallOfTheNasopharynx|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C111|PosteriorWallOfTheNasopharynx|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C111|PosteriorWallOfTheNasopharynx|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C111|PosteriorWallOfTheNasopharynx|808|LymphoepithelialCarcinoma|8085/3|SquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|808|LymphoepithelialCarcinoma|8086/3|SquamousCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C111|PosteriorWallOfTheNasopharynx|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C111|PosteriorWallOfTheNasopharynx|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C111|PosteriorWallOfTheNasopharynx|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C111|PosteriorWallOfTheNasopharynx|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C111|PosteriorWallOfTheNasopharynx|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C111|PosteriorWallOfTheNasopharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C111|PosteriorWallOfTheNasopharynx|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C111|PosteriorWallOfTheNasopharynx|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C111|PosteriorWallOfTheNasopharynx|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C111|PosteriorWallOfTheNasopharynx|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C111|PosteriorWallOfTheNasopharynx|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C111|PosteriorWallOfTheNasopharynx|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C111|PosteriorWallOfTheNasopharynx|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C111|PosteriorWallOfTheNasopharynx|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C111|PosteriorWallOfTheNasopharynx|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C111|PosteriorWallOfTheNasopharynx|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C111|PosteriorWallOfTheNasopharynx|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C111|PosteriorWallOfTheNasopharynx|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C111|PosteriorWallOfTheNasopharynx|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C111|PosteriorWallOfTheNasopharynx|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C111|PosteriorWallOfTheNasopharynx|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C111|PosteriorWallOfTheNasopharynx|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C111|PosteriorWallOfTheNasopharynx|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C111|PosteriorWallOfTheNasopharynx|872|Melanoma|8720/2|Stage0SkinMelanoma
C111|PosteriorWallOfTheNasopharynx|872|Melanoma|8720/3|Melanoma
C111|PosteriorWallOfTheNasopharynx|872|Melanoma|8721/3|NodularMelanoma
C111|PosteriorWallOfTheNasopharynx|872|Melanoma|8722/3|BalloonCellMelanoma
C111|PosteriorWallOfTheNasopharynx|872|Melanoma|8723/3|RegressingMelanoma
C111|PosteriorWallOfTheNasopharynx|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C111|PosteriorWallOfTheNasopharynx|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C111|PosteriorWallOfTheNasopharynx|874|Nevus|8745/3|DesmoplasticMelanoma
C111|PosteriorWallOfTheNasopharynx|874|Nevus|8746/3|MucosalLentiginousMelanoma
C111|PosteriorWallOfTheNasopharynx|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C111|PosteriorWallOfTheNasopharynx|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C111|PosteriorWallOfTheNasopharynx|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C111|PosteriorWallOfTheNasopharynx|880|Sarcoma|8800/3|Sarcoma
C111|PosteriorWallOfTheNasopharynx|880|Sarcoma|8801/3|SpindleCellSarcoma
C111|PosteriorWallOfTheNasopharynx|880|Sarcoma|8802/3|GiantCellSarcoma
C111|PosteriorWallOfTheNasopharynx|880|Sarcoma|8803/3|SmallCellSarcoma
C111|PosteriorWallOfTheNasopharynx|880|Sarcoma|8804/3|SarcomaEpithelioid
C111|PosteriorWallOfTheNasopharynx|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C111|PosteriorWallOfTheNasopharynx|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C111|PosteriorWallOfTheNasopharynx|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C111|PosteriorWallOfTheNasopharynx|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C111|PosteriorWallOfTheNasopharynx|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C111|PosteriorWallOfTheNasopharynx|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C111|PosteriorWallOfTheNasopharynx|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C111|PosteriorWallOfTheNasopharynx|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C111|PosteriorWallOfTheNasopharynx|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C111|PosteriorWallOfTheNasopharynx|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C111|PosteriorWallOfTheNasopharynx|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C111|PosteriorWallOfTheNasopharynx|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C111|PosteriorWallOfTheNasopharynx|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C111|PosteriorWallOfTheNasopharynx|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C111|PosteriorWallOfTheNasopharynx|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C111|PosteriorWallOfTheNasopharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C111|PosteriorWallOfTheNasopharynx|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C111|PosteriorWallOfTheNasopharynx|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C111|PosteriorWallOfTheNasopharynx|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C111|PosteriorWallOfTheNasopharynx|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C111|PosteriorWallOfTheNasopharynx|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C111|PosteriorWallOfTheNasopharynx|914|KaposiSarcoma|9140/3|KaposiSarcoma
C111|PosteriorWallOfTheNasopharynx|937|Chordoma|9370/3|Chordoma
C111|PosteriorWallOfTheNasopharynx|937|Chordoma|9371/3|ChondroidChordoma
C111|PosteriorWallOfTheNasopharynx|937|Chordoma|9372/3|DedifferentiatedChordoma
C111|PosteriorWallOfTheNasopharynx|959|Lymphoma|9590/3|Lymphoma
C111|PosteriorWallOfTheNasopharynx|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C111|PosteriorWallOfTheNasopharynx|959|Lymphoma|9596/3|CompositeLymphoma
C111|PosteriorWallOfTheNasopharynx|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C111|PosteriorWallOfTheNasopharynx|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C111|PosteriorWallOfTheNasopharynx|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C111|PosteriorWallOfTheNasopharynx|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C111|PosteriorWallOfTheNasopharynx|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C111|PosteriorWallOfTheNasopharynx|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C111|PosteriorWallOfTheNasopharynx|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C111|PosteriorWallOfTheNasopharynx|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C111|PosteriorWallOfTheNasopharynx|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C111|PosteriorWallOfTheNasopharynx|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C111|PosteriorWallOfTheNasopharynx|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C111|PosteriorWallOfTheNasopharynx|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C111|PosteriorWallOfTheNasopharynx|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C111|PosteriorWallOfTheNasopharynx|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C111|PosteriorWallOfTheNasopharynx|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C111|PosteriorWallOfTheNasopharynx|967|BCellLymphomas|9673/3|MantleCellLymphoma
C111|PosteriorWallOfTheNasopharynx|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C111|PosteriorWallOfTheNasopharynx|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C111|PosteriorWallOfTheNasopharynx|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C111|PosteriorWallOfTheNasopharynx|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C111|PosteriorWallOfTheNasopharynx|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C111|PosteriorWallOfTheNasopharynx|969|FollicularAdenoma|9690/3|LymphomaFollicular
C111|PosteriorWallOfTheNasopharynx|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C111|PosteriorWallOfTheNasopharynx|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C111|PosteriorWallOfTheNasopharynx|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C111|PosteriorWallOfTheNasopharynx|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C111|PosteriorWallOfTheNasopharynx|970|TCellLymphoma|9701/3|SezarySyndrome
C111|PosteriorWallOfTheNasopharynx|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C111|PosteriorWallOfTheNasopharynx|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C111|PosteriorWallOfTheNasopharynx|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C111|PosteriorWallOfTheNasopharynx|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C111|PosteriorWallOfTheNasopharynx|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C111|PosteriorWallOfTheNasopharynx|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C111|PosteriorWallOfTheNasopharynx|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C111|PosteriorWallOfTheNasopharynx|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C111|PosteriorWallOfTheNasopharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C111|PosteriorWallOfTheNasopharynx|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C111|PosteriorWallOfTheNasopharynx|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C111|PosteriorWallOfTheNasopharynx|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C111|PosteriorWallOfTheNasopharynx|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C111|PosteriorWallOfTheNasopharynx|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C111|PosteriorWallOfTheNasopharynx|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C111|PosteriorWallOfTheNasopharynx|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C111|PosteriorWallOfTheNasopharynx|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C111|PosteriorWallOfTheNasopharynx|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C111|PosteriorWallOfTheNasopharynx|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C111|PosteriorWallOfTheNasopharynx|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C111|PosteriorWallOfTheNasopharynx|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C111|PosteriorWallOfTheNasopharynx|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C111|PosteriorWallOfTheNasopharynx|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C111|PosteriorWallOfTheNasopharynx|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C111|PosteriorWallOfTheNasopharynx|981|PrecursorLymphoidNeoplasm|9812/3|null
C111|PosteriorWallOfTheNasopharynx|981|PrecursorLymphoidNeoplasm|9813/3|null
C111|PosteriorWallOfTheNasopharynx|981|PrecursorLymphoidNeoplasm|9814/3|null
C111|PosteriorWallOfTheNasopharynx|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C111|PosteriorWallOfTheNasopharynx|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C111|PosteriorWallOfTheNasopharynx|981|PrecursorLymphoidNeoplasm|9817/3|null
C111|PosteriorWallOfTheNasopharynx|981|PrecursorLymphoidNeoplasm|9818/3|null
C111|PosteriorWallOfTheNasopharynx|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C111|PosteriorWallOfTheNasopharynx|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C111|PosteriorWallOfTheNasopharynx|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C111|PosteriorWallOfTheNasopharynx|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C111|PosteriorWallOfTheNasopharynx|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C111|PosteriorWallOfTheNasopharynx|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C111|PosteriorWallOfTheNasopharynx|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8010/2|InSituCancer
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8010/3|CarcinomaNOSDNE
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8011/3|MalignantEpithelioma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8012/3|LargeCellCarcinoma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8014/3|LargeCellCarcinoma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8015/3|GlassyCellCarcinoma
C129-C132,C138-C139|Hypopharynx|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C129-C132,C138-C139|Hypopharynx|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C129-C132,C138-C139|Hypopharynx|802|Carcinoma|8022/3|PleomorphicCarcinoma
C129-C132,C138-C139|Hypopharynx|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C129-C132,C138-C139|Hypopharynx|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C129-C132,C138-C139|Hypopharynx|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C129-C132,C138-C139|Hypopharynx|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C129-C132,C138-C139|Hypopharynx|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C129-C132,C138-C139|Hypopharynx|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C129-C132,C138-C139|Hypopharynx|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C129-C132,C138-C139|Hypopharynx|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C129-C132,C138-C139|Hypopharynx|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C129-C132,C138-C139|Hypopharynx|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C129-C132,C138-C139|Hypopharynx|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C129-C132,C138-C139|Hypopharynx|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C129-C132,C138-C139|Hypopharynx|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C129-C132,C138-C139|Hypopharynx|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C129-C132,C138-C139|Hypopharynx|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C129-C132,C138-C139|Hypopharynx|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C129-C132,C138-C139|Hypopharynx|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C129-C132,C138-C139|Hypopharynx|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C129-C132,C138-C139|Hypopharynx|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C129-C132,C138-C139|Hypopharynx|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C129-C132,C138-C139|Hypopharynx|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C129-C132,C138-C139|Hypopharynx|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C129-C132,C138-C139|Hypopharynx|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C129-C132,C138-C139|Hypopharynx|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C129-C132,C138-C139|Hypopharynx|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C129-C132,C138-C139|Hypopharynx|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C129-C132,C138-C139|Hypopharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C129-C132,C138-C139|Hypopharynx|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C129-C132,C138-C139|Hypopharynx|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C129-C132,C138-C139|Hypopharynx|914|KaposiSarcoma|9140/3|KaposiSarcoma
C129-C132,C138-C139|Hypopharynx|959|Lymphoma|9590/3|Lymphoma
C129-C132,C138-C139|Hypopharynx|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C129-C132,C138-C139|Hypopharynx|959|Lymphoma|9596/3|CompositeLymphoma
C129-C132,C138-C139|Hypopharynx|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C129-C132,C138-C139|Hypopharynx|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C129-C132,C138-C139|Hypopharynx|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C129-C132,C138-C139|Hypopharynx|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C129-C132,C138-C139|Hypopharynx|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C129-C132,C138-C139|Hypopharynx|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C129-C132,C138-C139|Hypopharynx|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C129-C132,C138-C139|Hypopharynx|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C129-C132,C138-C139|Hypopharynx|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C129-C132,C138-C139|Hypopharynx|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C129-C132,C138-C139|Hypopharynx|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C129-C132,C138-C139|Hypopharynx|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C129-C132,C138-C139|Hypopharynx|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C129-C132,C138-C139|Hypopharynx|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C129-C132,C138-C139|Hypopharynx|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C129-C132,C138-C139|Hypopharynx|967|BCellLymphomas|9673/3|MantleCellLymphoma
C129-C132,C138-C139|Hypopharynx|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C129-C132,C138-C139|Hypopharynx|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C129-C132,C138-C139|Hypopharynx|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C129-C132,C138-C139|Hypopharynx|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C129-C132,C138-C139|Hypopharynx|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C129-C132,C138-C139|Hypopharynx|969|FollicularAdenoma|9690/3|LymphomaFollicular
C129-C132,C138-C139|Hypopharynx|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C129-C132,C138-C139|Hypopharynx|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C129-C132,C138-C139|Hypopharynx|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C129-C132,C138-C139|Hypopharynx|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C129-C132,C138-C139|Hypopharynx|970|TCellLymphoma|9701/3|SezarySyndrome
C129-C132,C138-C139|Hypopharynx|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C129-C132,C138-C139|Hypopharynx|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C129-C132,C138-C139|Hypopharynx|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C129-C132,C138-C139|Hypopharynx|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C129-C132,C138-C139|Hypopharynx|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C129-C132,C138-C139|Hypopharynx|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C129-C132,C138-C139|Hypopharynx|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C129-C132,C138-C139|Hypopharynx|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C129-C132,C138-C139|Hypopharynx|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C129-C132,C138-C139|Hypopharynx|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C129-C132,C138-C139|Hypopharynx|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C129-C132,C138-C139|Hypopharynx|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C129-C132,C138-C139|Hypopharynx|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C129-C132,C138-C139|Hypopharynx|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C129-C132,C138-C139|Hypopharynx|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C129-C132,C138-C139|Hypopharynx|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C129-C132,C138-C139|Hypopharynx|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C129-C132,C138-C139|Hypopharynx|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C129-C132,C138-C139|Hypopharynx|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C129-C132,C138-C139|Hypopharynx|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C129-C132,C138-C139|Hypopharynx|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C129-C132,C138-C139|Hypopharynx|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9812/3|null
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9813/3|null
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9814/3|null
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9817/3|null
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9818/3|null
C129-C132,C138-C139|Hypopharynx|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C129-C132,C138-C139|Hypopharynx|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C129-C132,C138-C139|Hypopharynx|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C129-C132,C138-C139|Hypopharynx|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C129-C132,C138-C139|Hypopharynx|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C129-C132,C138-C139|Hypopharynx|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C129-C132,C138-C139|Hypopharynx|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C129-C132,C138-C139|Hypopharynx|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C140,C142,C148|Pharynx|801|Carcinoma|8010/2|InSituCancer
C140,C142,C148|Pharynx|801|Carcinoma|8010/3|CarcinomaNOSDNE
C140,C142,C148|Pharynx|801|Carcinoma|8011/3|MalignantEpithelioma
C140,C142,C148|Pharynx|801|Carcinoma|8012/3|LargeCellCarcinoma
C140,C142,C148|Pharynx|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C140,C142,C148|Pharynx|801|Carcinoma|8014/3|LargeCellCarcinoma
C140,C142,C148|Pharynx|801|Carcinoma|8015/3|GlassyCellCarcinoma
C140,C142,C148|Pharynx|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C140,C142,C148|Pharynx|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C140,C142,C148|Pharynx|802|Carcinoma|8022/3|PleomorphicCarcinoma
C140,C142,C148|Pharynx|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C140,C142,C148|Pharynx|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C140,C142,C148|Pharynx|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C140,C142,C148|Pharynx|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C140,C142,C148|Pharynx|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C140,C142,C148|Pharynx|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C140,C142,C148|Pharynx|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C140,C142,C148|Pharynx|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C140,C142,C148|Pharynx|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C140,C142,C148|Pharynx|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C140,C142,C148|Pharynx|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C140,C142,C148|Pharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C140,C142,C148|Pharynx|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C140,C142,C148|Pharynx|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C140,C142,C148|Pharynx|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C140,C142,C148|Pharynx|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C140,C142,C148|Pharynx|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C140,C142,C148|Pharynx|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C140,C142,C148|Pharynx|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C140,C142,C148|Pharynx|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C140,C142,C148|Pharynx|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C140,C142,C148|Pharynx|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C140,C142,C148|Pharynx|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C140,C142,C148|Pharynx|889|MyomatousNeoplasm|8895/3|Myosarcoma
C140,C142,C148|Pharynx|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C140,C142,C148|Pharynx|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C140,C142,C148|Pharynx|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C140,C142,C148|Pharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C140,C142,C148|Pharynx|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C140,C142,C148|Pharynx|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C140,C142,C148|Pharynx|937|Chordoma|9370/3|Chordoma
C140,C142,C148|Pharynx|937|Chordoma|9371/3|ChondroidChordoma
C140,C142,C148|Pharynx|937|Chordoma|9372/3|DedifferentiatedChordoma
C140,C142,C148|Pharynx|959|Lymphoma|9590/3|Lymphoma
C140,C142,C148|Pharynx|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C140,C142,C148|Pharynx|959|Lymphoma|9596/3|CompositeLymphoma
C140,C142,C148|Pharynx|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C140,C142,C148|Pharynx|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C140,C142,C148|Pharynx|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C140,C142,C148|Pharynx|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C140,C142,C148|Pharynx|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C140,C142,C148|Pharynx|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C140,C142,C148|Pharynx|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C140,C142,C148|Pharynx|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C140,C142,C148|Pharynx|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C140,C142,C148|Pharynx|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C140,C142,C148|Pharynx|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C140,C142,C148|Pharynx|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C140,C142,C148|Pharynx|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C140,C142,C148|Pharynx|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C140,C142,C148|Pharynx|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C140,C142,C148|Pharynx|967|BCellLymphomas|9673/3|MantleCellLymphoma
C140,C142,C148|Pharynx|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C140,C142,C148|Pharynx|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C140,C142,C148|Pharynx|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C140,C142,C148|Pharynx|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C140,C142,C148|Pharynx|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C140,C142,C148|Pharynx|969|FollicularAdenoma|9690/3|LymphomaFollicular
C140,C142,C148|Pharynx|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C140,C142,C148|Pharynx|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C140,C142,C148|Pharynx|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C140,C142,C148|Pharynx|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C140,C142,C148|Pharynx|970|TCellLymphoma|9701/3|SezarySyndrome
C140,C142,C148|Pharynx|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C140,C142,C148|Pharynx|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C140,C142,C148|Pharynx|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C140,C142,C148|Pharynx|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C140,C142,C148|Pharynx|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C140,C142,C148|Pharynx|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C140,C142,C148|Pharynx|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C140,C142,C148|Pharynx|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C140,C142,C148|Pharynx|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C140,C142,C148|Pharynx|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C140,C142,C148|Pharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C140,C142,C148|Pharynx|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C140,C142,C148|Pharynx|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C140,C142,C148|Pharynx|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C140,C142,C148|Pharynx|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C140,C142,C148|Pharynx|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C140,C142,C148|Pharynx|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C140,C142,C148|Pharynx|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C140,C142,C148|Pharynx|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C140,C142,C148|Pharynx|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C140,C142,C148|Pharynx|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C140,C142,C148|Pharynx|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C140,C142,C148|Pharynx|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9812/3|null
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9813/3|null
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9814/3|null
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9817/3|null
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9818/3|null
C140,C142,C148|Pharynx|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C140,C142,C148|Pharynx|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C140,C142,C148|Pharynx|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C140,C142,C148|Pharynx|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C140,C142,C148|Pharynx|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C140,C142,C148|Pharynx|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C140,C142,C148|Pharynx|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C140,C142,C148|Pharynx|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C150-C155,C158-C159|Esophagus|801|Carcinoma|8010/2|InSituCancer
C150-C155,C158-C159|Esophagus|801|Carcinoma|8010/3|CarcinomaNOSDNE
C150-C155,C158-C159|Esophagus|801|Carcinoma|8011/3|MalignantEpithelioma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8012/3|LargeCellCarcinoma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8014/3|LargeCellCarcinoma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8015/3|GlassyCellCarcinoma
C150-C155,C158-C159|Esophagus|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C150-C155,C158-C159|Esophagus|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C150-C155,C158-C159|Esophagus|802|Carcinoma|8022/3|PleomorphicCarcinoma
C150-C155,C158-C159|Esophagus|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C150-C155,C158-C159|Esophagus|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C150-C155,C158-C159|Esophagus|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C150-C155,C158-C159|Esophagus|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C150-C155,C158-C159|Esophagus|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C150-C155,C158-C159|Esophagus|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C150-C155,C158-C159|Esophagus|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C150-C155,C158-C159|Esophagus|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C150-C155,C158-C159|Esophagus|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C150-C155,C158-C159|Esophagus|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C150-C155,C158-C159|Esophagus|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C150-C155,C158-C159|Esophagus|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C150-C155,C158-C159|Esophagus|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8145/3|DiffuseTypeAdenocarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C150-C155,C158-C159|Esophagus|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C150-C155,C158-C159|Esophagus|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C150-C155,C158-C159|Esophagus|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C150-C155,C158-C159|Esophagus|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C150-C155,C158-C159|Esophagus|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C150-C155,C158-C159|Esophagus|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C150-C155,C158-C159|Esophagus|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C150-C155,C158-C159|Esophagus|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C150-C155,C158-C159|Esophagus|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C150-C155,C158-C159|Esophagus|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C150-C155,C158-C159|Esophagus|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C150-C155,C158-C159|Esophagus|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C150-C155,C158-C159|Esophagus|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C150-C155,C158-C159|Esophagus|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C150-C155,C158-C159|Esophagus|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C150-C155,C158-C159|Esophagus|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C150-C155,C158-C159|Esophagus|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C150-C155,C158-C159|Esophagus|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C150-C155,C158-C159|Esophagus|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C150-C155,C158-C159|Esophagus|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C150-C155,C158-C159|Esophagus|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C150-C155,C158-C159|Esophagus|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C150-C155,C158-C159|Esophagus|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C150-C155,C158-C159|Esophagus|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C150-C155,C158-C159|Esophagus|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8720/2|Stage0SkinMelanoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8720/3|Melanoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8721/3|NodularMelanoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8722/3|BalloonCellMelanoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8723/3|RegressingMelanoma
C150-C155,C158-C159|Esophagus|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C150-C155,C158-C159|Esophagus|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C150-C155,C158-C159|Esophagus|874|Nevus|8745/3|DesmoplasticMelanoma
C150-C155,C158-C159|Esophagus|874|Nevus|8746/3|MucosalLentiginousMelanoma
C150-C155,C158-C159|Esophagus|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C150-C155,C158-C159|Esophagus|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C150-C155,C158-C159|Esophagus|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C150-C155,C158-C159|Esophagus|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C150-C155,C158-C159|Esophagus|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C150-C155,C158-C159|Esophagus|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C150-C155,C158-C159|Esophagus|889|MyomatousNeoplasm|8895/3|Myosarcoma
C150-C155,C158-C159|Esophagus|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C150-C155,C158-C159|Esophagus|898|Carcinosarcoma|8980/3|Carcinosarcoma
C150-C155,C158-C159|Esophagus|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C150-C155,C158-C159|Esophagus|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C150-C155,C158-C159|Esophagus|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C150-C155,C158-C159|Esophagus|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C150-C155,C158-C159|Esophagus|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C150-C155,C158-C159|Esophagus|970|TCellLymphoma|9701/3|SezarySyndrome
C150-C155,C158-C159|Esophagus|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C150-C155,C158-C159|Esophagus|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C150-C155,C158-C159|Esophagus|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C150-C155,C158-C159|Esophagus|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C150-C155,C158-C159|Esophagus|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C150-C155,C158-C159|Esophagus|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C150-C155,C158-C159|Esophagus|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C150-C155,C158-C159|Esophagus|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C150-C155,C158-C159|Esophagus|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C150-C155,C158-C159|Esophagus|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9731/3|Plasmacytoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C150-C155,C158-C159|Esophagus|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C150-C155,C158-C159|Esophagus|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C150-C155,C158-C159|Esophagus|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C150-C155,C158-C159|Esophagus|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C150-C155,C158-C159|Esophagus|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C150-C155,C158-C159|Esophagus|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C150-C155,C158-C159|Esophagus|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C150-C155,C158-C159|Esophagus|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C150-C155,C158-C159|Esophagus|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C150-C155,C158-C159|Esophagus|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C150-C155,C158-C159|Esophagus|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C150-C155,C158-C159|Esophagus|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9812/3|null
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9813/3|null
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9814/3|null
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9817/3|null
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9818/3|null
C150-C155,C158-C159|Esophagus|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C150-C155,C158-C159|Esophagus|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C150-C155,C158-C159|Esophagus|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C150-C155,C158-C159|Esophagus|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C150-C155,C158-C159|Esophagus|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C150-C155,C158-C159|Esophagus|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C150-C155,C158-C159|Esophagus|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C150-C155,C158-C159|Esophagus|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C160-C166,C168-C169|Stomach|801|Carcinoma|8010/2|InSituCancer
C160-C166,C168-C169|Stomach|801|Carcinoma|8010/3|CarcinomaNOSDNE
C160-C166,C168-C169|Stomach|801|Carcinoma|8011/3|MalignantEpithelioma
C160-C166,C168-C169|Stomach|801|Carcinoma|8012/3|LargeCellCarcinoma
C160-C166,C168-C169|Stomach|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C160-C166,C168-C169|Stomach|801|Carcinoma|8014/3|LargeCellCarcinoma
C160-C166,C168-C169|Stomach|801|Carcinoma|8015/3|GlassyCellCarcinoma
C160-C166,C168-C169|Stomach|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C160-C166,C168-C169|Stomach|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C160-C166,C168-C169|Stomach|802|Carcinoma|8022/3|PleomorphicCarcinoma
C160-C166,C168-C169|Stomach|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C160-C166,C168-C169|Stomach|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C160-C166,C168-C169|Stomach|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C160-C166,C168-C169|Stomach|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C160-C166,C168-C169|Stomach|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C160-C166,C168-C169|Stomach|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C160-C166,C168-C169|Stomach|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C160-C166,C168-C169|Stomach|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C160-C166,C168-C169|Stomach|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C160-C166,C168-C169|Stomach|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C160-C166,C168-C169|Stomach|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C160-C166,C168-C169|Stomach|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C160-C166,C168-C169|Stomach|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C160-C166,C168-C169|Stomach|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C160-C166,C168-C169|Stomach|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8140/3|Adenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8142/3|LinitisPlastica
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8144/3|IntestinalTypeAdenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8145/3|DiffuseTypeAdenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C160-C166,C168-C169|Stomach|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C160-C166,C168-C169|Stomach|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C160-C166,C168-C169|Stomach|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C160-C166,C168-C169|Stomach|821|AdenocarcinomaInAdenomatousPolyp|8214/3|GastricParietalCellAdenocarcinoma
C160-C166,C168-C169|Stomach|822|FamilialAdenomatousPolyposis|8220/2|AdenocarcinomaInSitu
C160-C166,C168-C169|Stomach|822|FamilialAdenomatousPolyposis|8220/3|FamilialAdenomatousPolyposis
C160-C166,C168-C169|Stomach|822|FamilialAdenomatousPolyposis|8221/2|AdenomatousPolyp
C160-C166,C168-C169|Stomach|822|FamilialAdenomatousPolyposis|8221/3|AdenomatousPolyp
C160-C166,C168-C169|Stomach|823|SolidCarcinoma|8230/2|InSituCancer
C160-C166,C168-C169|Stomach|823|SolidCarcinoma|8230/3|SolidCarcinoma
C160-C166,C168-C169|Stomach|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C160-C166,C168-C169|Stomach|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C160-C166,C168-C169|Stomach|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C160-C166,C168-C169|Stomach|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C160-C166,C168-C169|Stomach|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C160-C166,C168-C169|Stomach|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C160-C166,C168-C169|Stomach|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C160-C166,C168-C169|Stomach|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C160-C166,C168-C169|Stomach|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C160-C166,C168-C169|Stomach|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C160-C166,C168-C169|Stomach|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C160-C166,C168-C169|Stomach|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C160-C166,C168-C169|Stomach|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C160-C166,C168-C169|Stomach|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C160-C166,C168-C169|Stomach|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C160-C166,C168-C169|Stomach|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C160-C166,C168-C169|Stomach|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C160-C166,C168-C169|Stomach|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C160-C166,C168-C169|Stomach|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C160-C166,C168-C169|Stomach|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C160-C166,C168-C169|Stomach|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C160-C166,C168-C169|Stomach|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C160-C166,C168-C169|Stomach|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C160-C166,C168-C169|Stomach|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C160-C166,C168-C169|Stomach|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C160-C166,C168-C169|Stomach|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C160-C166,C168-C169|Stomach|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C160-C166,C168-C169|Stomach|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C160-C166,C168-C169|Stomach|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C160-C166,C168-C169|Stomach|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8800/3|Sarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8801/3|SpindleCellSarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8802/3|GiantCellSarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8803/3|SmallCellSarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8804/3|SarcomaEpithelioid
C160-C166,C168-C169|Stomach|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C160-C166,C168-C169|Stomach|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C160-C166,C168-C169|Stomach|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C160-C166,C168-C169|Stomach|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C160-C166,C168-C169|Stomach|889|MyomatousNeoplasm|8895/3|Myosarcoma
C160-C166,C168-C169|Stomach|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C160-C166,C168-C169|Stomach|893|StromalSarcoma|8934/3|Carcinofibroma
C160-C166,C168-C169|Stomach|893|StromalSarcoma|8935/3|StromalSarcoma
C160-C166,C168-C169|Stomach|893|StromalSarcoma|8936/3|HighRiskGastrointestinalStromalTumor
C160-C166,C168-C169|Stomach|898|Carcinosarcoma|8980/3|Carcinosarcoma
C160-C166,C168-C169|Stomach|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C160-C166,C168-C169|Stomach|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C160-C166,C168-C169|Stomach|959|Lymphoma|9590/3|Lymphoma
C160-C166,C168-C169|Stomach|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C160-C166,C168-C169|Stomach|959|Lymphoma|9596/3|CompositeLymphoma
C160-C166,C168-C169|Stomach|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C160-C166,C168-C169|Stomach|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C160-C166,C168-C169|Stomach|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C160-C166,C168-C169|Stomach|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C160-C166,C168-C169|Stomach|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C160-C166,C168-C169|Stomach|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C160-C166,C168-C169|Stomach|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C160-C166,C168-C169|Stomach|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C160-C166,C168-C169|Stomach|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C160-C166,C168-C169|Stomach|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C160-C166,C168-C169|Stomach|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C160-C166,C168-C169|Stomach|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C160-C166,C168-C169|Stomach|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C160-C166,C168-C169|Stomach|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C160-C166,C168-C169|Stomach|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C160-C166,C168-C169|Stomach|967|BCellLymphomas|9673/3|MantleCellLymphoma
C160-C166,C168-C169|Stomach|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C160-C166,C168-C169|Stomach|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C160-C166,C168-C169|Stomach|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C160-C166,C168-C169|Stomach|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C160-C166,C168-C169|Stomach|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C160-C166,C168-C169|Stomach|969|FollicularAdenoma|9690/3|LymphomaFollicular
C160-C166,C168-C169|Stomach|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C160-C166,C168-C169|Stomach|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C160-C166,C168-C169|Stomach|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C160-C166,C168-C169|Stomach|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C160-C166,C168-C169|Stomach|970|TCellLymphoma|9701/3|SezarySyndrome
C160-C166,C168-C169|Stomach|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C160-C166,C168-C169|Stomach|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C160-C166,C168-C169|Stomach|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C160-C166,C168-C169|Stomach|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C160-C166,C168-C169|Stomach|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C160-C166,C168-C169|Stomach|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C160-C166,C168-C169|Stomach|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C160-C166,C168-C169|Stomach|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C160-C166,C168-C169|Stomach|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C160-C166,C168-C169|Stomach|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9731/3|Plasmacytoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9732/3|PlasmaCellMyeloma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C160-C166,C168-C169|Stomach|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C160-C166,C168-C169|Stomach|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C160-C166,C168-C169|Stomach|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C160-C166,C168-C169|Stomach|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C160-C166,C168-C169|Stomach|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C160-C166,C168-C169|Stomach|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C160-C166,C168-C169|Stomach|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C160-C166,C168-C169|Stomach|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C160-C166,C168-C169|Stomach|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C160-C166,C168-C169|Stomach|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C160-C166,C168-C169|Stomach|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C160-C166,C168-C169|Stomach|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9812/3|null
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9813/3|null
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9814/3|null
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9817/3|null
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9818/3|null
C160-C166,C168-C169|Stomach|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C160-C166,C168-C169|Stomach|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C160-C166,C168-C169|Stomach|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C160-C166,C168-C169|Stomach|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C160-C166,C168-C169|Stomach|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C160-C166,C168-C169|Stomach|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C160-C166,C168-C169|Stomach|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C160-C166,C168-C169|Stomach|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C170-C173,C178-C179|SmallIntestine|801|Carcinoma|8010/2|InSituCancer
C170-C173,C178-C179|SmallIntestine|801|Carcinoma|8010/3|CarcinomaNOSDNE
C170-C173,C178-C179|SmallIntestine|801|Carcinoma|8011/3|MalignantEpithelioma
C170-C173,C178-C179|SmallIntestine|801|Carcinoma|8012/3|LargeCellCarcinoma
C170-C173,C178-C179|SmallIntestine|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C170-C173,C178-C179|SmallIntestine|801|Carcinoma|8014/3|LargeCellCarcinoma
C170-C173,C178-C179|SmallIntestine|801|Carcinoma|8015/3|GlassyCellCarcinoma
C170-C173,C178-C179|SmallIntestine|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C170-C173,C178-C179|SmallIntestine|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C170-C173,C178-C179|SmallIntestine|802|Carcinoma|8022/3|PleomorphicCarcinoma
C170-C173,C178-C179|SmallIntestine|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C170-C173,C178-C179|SmallIntestine|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C170-C173,C178-C179|SmallIntestine|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C170-C173,C178-C179|SmallIntestine|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C170-C173,C178-C179|SmallIntestine|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C170-C173,C178-C179|SmallIntestine|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C170-C173,C178-C179|SmallIntestine|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C170-C173,C178-C179|SmallIntestine|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C170-C173,C178-C179|SmallIntestine|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C170-C173,C178-C179|SmallIntestine|814|Adenocarcinoma|8140/3|Adenocarcinoma
C170-C173,C178-C179|SmallIntestine|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C170-C173,C178-C179|SmallIntestine|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C170-C173,C178-C179|SmallIntestine|814|Adenocarcinoma|8145/3|DiffuseTypeAdenocarcinoma
C170-C173,C178-C179|SmallIntestine|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C170-C173,C178-C179|SmallIntestine|815|EndocrineGlandNeoplasms|8152/3|MalignantPancreaticGlucagonoma
C170-C173,C178-C179|SmallIntestine|815|EndocrineGlandNeoplasms|8153/3|MalignantGastrinoma
C170-C173,C178-C179|SmallIntestine|815|EndocrineGlandNeoplasms|8156/3|MalignantSomatostatinoma
C170-C173,C178-C179|SmallIntestine|815|EndocrineGlandNeoplasms|8157/3|MalignantEnteroglucagonoma
C170-C173,C178-C179|SmallIntestine|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C170-C173,C178-C179|SmallIntestine|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C170-C173,C178-C179|SmallIntestine|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C170-C173,C178-C179|SmallIntestine|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C170-C173,C178-C179|SmallIntestine|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C170-C173,C178-C179|SmallIntestine|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C170-C173,C178-C179|SmallIntestine|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C170-C173,C178-C179|SmallIntestine|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C170-C173,C178-C179|SmallIntestine|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C170-C173,C178-C179|SmallIntestine|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C170-C173,C178-C179|SmallIntestine|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C170-C173,C178-C179|SmallIntestine|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C170-C173,C178-C179|SmallIntestine|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C170-C173,C178-C179|SmallIntestine|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C170-C173,C178-C179|SmallIntestine|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C170-C173,C178-C179|SmallIntestine|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C170-C173,C178-C179|SmallIntestine|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C170-C173,C178-C179|SmallIntestine|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C170-C173,C178-C179|SmallIntestine|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C170-C173,C178-C179|SmallIntestine|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C170-C173,C178-C179|SmallIntestine|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C170-C173,C178-C179|SmallIntestine|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C170-C173,C178-C179|SmallIntestine|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C170-C173,C178-C179|SmallIntestine|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C170-C173,C178-C179|SmallIntestine|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C170-C173,C178-C179|SmallIntestine|871|MalignantGlomusTumor|8710/3|MalignantGlomusTumor
C170-C173,C178-C179|SmallIntestine|880|Sarcoma|8800/3|Sarcoma
C170-C173,C178-C179|SmallIntestine|880|Sarcoma|8801/3|SpindleCellSarcoma
C170-C173,C178-C179|SmallIntestine|880|Sarcoma|8802/3|GiantCellSarcoma
C170-C173,C178-C179|SmallIntestine|880|Sarcoma|8803/3|SmallCellSarcoma
C170-C173,C178-C179|SmallIntestine|880|Sarcoma|8804/3|SarcomaEpithelioid
C170-C173,C178-C179|SmallIntestine|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C170-C173,C178-C179|SmallIntestine|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C170-C173,C178-C179|SmallIntestine|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C170-C173,C178-C179|SmallIntestine|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C170-C173,C178-C179|SmallIntestine|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C170-C173,C178-C179|SmallIntestine|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C170-C173,C178-C179|SmallIntestine|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C170-C173,C178-C179|SmallIntestine|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C170-C173,C178-C179|SmallIntestine|885|Liposarcoma|8850/3|Liposarcoma
C170-C173,C178-C179|SmallIntestine|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C170-C173,C178-C179|SmallIntestine|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C170-C173,C178-C179|SmallIntestine|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C170-C173,C178-C179|SmallIntestine|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C170-C173,C178-C179|SmallIntestine|885|Liposarcoma|8855/3|Liposarcoma
C170-C173,C178-C179|SmallIntestine|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C170-C173,C178-C179|SmallIntestine|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C170-C173,C178-C179|SmallIntestine|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C170-C173,C178-C179|SmallIntestine|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C170-C173,C178-C179|SmallIntestine|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C170-C173,C178-C179|SmallIntestine|889|MyomatousNeoplasm|8895/3|Myosarcoma
C170-C173,C178-C179|SmallIntestine|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C170-C173,C178-C179|SmallIntestine|893|StromalSarcoma|8934/3|Carcinofibroma
C170-C173,C178-C179|SmallIntestine|893|StromalSarcoma|8935/3|StromalSarcoma
C170-C173,C178-C179|SmallIntestine|893|StromalSarcoma|8936/3|HighRiskGastrointestinalStromalTumor
C170-C173,C178-C179|SmallIntestine|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C170-C173,C178-C179|SmallIntestine|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C170-C173,C178-C179|SmallIntestine|959|Lymphoma|9590/3|Lymphoma
C170-C173,C178-C179|SmallIntestine|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C170-C173,C178-C179|SmallIntestine|959|Lymphoma|9596/3|CompositeLymphoma
C170-C173,C178-C179|SmallIntestine|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C170-C173,C178-C179|SmallIntestine|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C170-C173,C178-C179|SmallIntestine|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C170-C173,C178-C179|SmallIntestine|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C170-C173,C178-C179|SmallIntestine|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C170-C173,C178-C179|SmallIntestine|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C170-C173,C178-C179|SmallIntestine|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C170-C173,C178-C179|SmallIntestine|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C170-C173,C178-C179|SmallIntestine|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C170-C173,C178-C179|SmallIntestine|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C170-C173,C178-C179|SmallIntestine|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C170-C173,C178-C179|SmallIntestine|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C170-C173,C178-C179|SmallIntestine|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C170-C173,C178-C179|SmallIntestine|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C170-C173,C178-C179|SmallIntestine|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C170-C173,C178-C179|SmallIntestine|967|BCellLymphomas|9673/3|MantleCellLymphoma
C170-C173,C178-C179|SmallIntestine|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C170-C173,C178-C179|SmallIntestine|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C170-C173,C178-C179|SmallIntestine|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C170-C173,C178-C179|SmallIntestine|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C170-C173,C178-C179|SmallIntestine|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C170-C173,C178-C179|SmallIntestine|969|FollicularAdenoma|9690/3|LymphomaFollicular
C170-C173,C178-C179|SmallIntestine|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C170-C173,C178-C179|SmallIntestine|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C170-C173,C178-C179|SmallIntestine|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C170-C173,C178-C179|SmallIntestine|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C170-C173,C178-C179|SmallIntestine|970|TCellLymphoma|9701/3|SezarySyndrome
C170-C173,C178-C179|SmallIntestine|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C170-C173,C178-C179|SmallIntestine|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C170-C173,C178-C179|SmallIntestine|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C170-C173,C178-C179|SmallIntestine|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C170-C173,C178-C179|SmallIntestine|971|AdultNonHodgkinLymphoma|9717/3|IntestinalTCellLymphomaNOS
C170-C173,C178-C179|SmallIntestine|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C170-C173,C178-C179|SmallIntestine|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C170-C173,C178-C179|SmallIntestine|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C170-C173,C178-C179|SmallIntestine|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C170-C173,C178-C179|SmallIntestine|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C170-C173,C178-C179|SmallIntestine|973|Plasmacytoma|9731/3|Plasmacytoma
C170-C173,C178-C179|SmallIntestine|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C170-C173,C178-C179|SmallIntestine|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C170-C173,C178-C179|SmallIntestine|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C170-C173,C178-C179|SmallIntestine|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C170-C173,C178-C179|SmallIntestine|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C170-C173,C178-C179|SmallIntestine|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C170-C173,C178-C179|SmallIntestine|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C170-C173,C178-C179|SmallIntestine|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C170-C173,C178-C179|SmallIntestine|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C170-C173,C178-C179|SmallIntestine|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C170-C173,C178-C179|SmallIntestine|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C170-C173,C178-C179|SmallIntestine|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C170-C173,C178-C179|SmallIntestine|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C170-C173,C178-C179|SmallIntestine|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C170-C173,C178-C179|SmallIntestine|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C170-C173,C178-C179|SmallIntestine|976|ImmunoproliferativeDisorder|9764/3|ImmunoproliferativeDisorder
C170-C173,C178-C179|SmallIntestine|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9812/3|null
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9813/3|null
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9814/3|null
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9817/3|null
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9818/3|null
C170-C173,C178-C179|SmallIntestine|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C170-C173,C178-C179|SmallIntestine|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C170-C173,C178-C179|SmallIntestine|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C170-C173,C178-C179|SmallIntestine|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C170-C173,C178-C179|SmallIntestine|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C170-C173,C178-C179|SmallIntestine|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C170-C173,C178-C179|SmallIntestine|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C170-C173,C178-C179|SmallIntestine|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C180, C182-C189, C199|LargeIntestine|801|Carcinoma|8010/2|InSituCancer
C180, C182-C189, C199|LargeIntestine|801|Carcinoma|8010/3|CarcinomaNOSDNE
C180, C182-C189, C199|LargeIntestine|801|Carcinoma|8011/3|MalignantEpithelioma
C180, C182-C189, C199|LargeIntestine|801|Carcinoma|8012/3|LargeCellCarcinoma
C180, C182-C189, C199|LargeIntestine|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C180, C182-C189, C199|LargeIntestine|801|Carcinoma|8014/3|LargeCellCarcinoma
C180, C182-C189, C199|LargeIntestine|801|Carcinoma|8015/3|GlassyCellCarcinoma
C180, C182-C189, C199|LargeIntestine|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C180, C182-C189, C199|LargeIntestine|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C180, C182-C189, C199|LargeIntestine|802|Carcinoma|8022/3|PleomorphicCarcinoma
C180, C182-C189, C199|LargeIntestine|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C180, C182-C189, C199|LargeIntestine|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C180, C182-C189, C199|LargeIntestine|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C180, C182-C189, C199|LargeIntestine|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C180, C182-C189, C199|LargeIntestine|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C180, C182-C189, C199|LargeIntestine|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C180, C182-C189, C199|LargeIntestine|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C180, C182-C189, C199|LargeIntestine|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C180, C182-C189, C199|LargeIntestine|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C180, C182-C189, C199|LargeIntestine|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C180, C182-C189, C199|LargeIntestine|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C180, C182-C189, C199|LargeIntestine|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C180, C182-C189, C199|LargeIntestine|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C180, C182-C189, C199|LargeIntestine|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C180, C182-C189, C199|LargeIntestine|814|Adenocarcinoma|8140/3|Adenocarcinoma
C180, C182-C189, C199|LargeIntestine|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|814|Adenocarcinoma|8145/3|DiffuseTypeAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C180, C182-C189, C199|LargeIntestine|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C180, C182-C189, C199|LargeIntestine|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C180, C182-C189, C199|LargeIntestine|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|821|AdenocarcinomaInAdenomatousPolyp|8213/3|SerratedAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|822|FamilialAdenomatousPolyposis|8220/2|AdenocarcinomaInSitu
C180, C182-C189, C199|LargeIntestine|822|FamilialAdenomatousPolyposis|8220/3|FamilialAdenomatousPolyposis
C180, C182-C189, C199|LargeIntestine|822|FamilialAdenomatousPolyposis|8221/2|AdenomatousPolyp
C180, C182-C189, C199|LargeIntestine|822|FamilialAdenomatousPolyposis|8221/3|AdenomatousPolyp
C180, C182-C189, C199|LargeIntestine|823|SolidCarcinoma|8230/2|InSituCancer
C180, C182-C189, C199|LargeIntestine|823|SolidCarcinoma|8230/3|SolidCarcinoma
C180, C182-C189, C199|LargeIntestine|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C180, C182-C189, C199|LargeIntestine|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C180, C182-C189, C199|LargeIntestine|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C180, C182-C189, C199|LargeIntestine|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C180, C182-C189, C199|LargeIntestine|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C180, C182-C189, C199|LargeIntestine|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C180, C182-C189, C199|LargeIntestine|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C180, C182-C189, C199|LargeIntestine|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C180, C182-C189, C199|LargeIntestine|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C180, C182-C189, C199|LargeIntestine|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C180, C182-C189, C199|LargeIntestine|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C180, C182-C189, C199|LargeIntestine|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C180, C182-C189, C199|LargeIntestine|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C180, C182-C189, C199|LargeIntestine|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C180, C182-C189, C199|LargeIntestine|826|PapillaryAdenocarcinoma|8265/3|MicropapillaryCarcinoma
C180, C182-C189, C199|LargeIntestine|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C180, C182-C189, C199|LargeIntestine|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C180, C182-C189, C199|LargeIntestine|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C180, C182-C189, C199|LargeIntestine|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C180, C182-C189, C199|LargeIntestine|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C180, C182-C189, C199|LargeIntestine|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C180, C182-C189, C199|LargeIntestine|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C180, C182-C189, C199|LargeIntestine|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C180, C182-C189, C199|LargeIntestine|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C180, C182-C189, C199|LargeIntestine|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C180, C182-C189, C199|LargeIntestine|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C180, C182-C189, C199|LargeIntestine|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C180, C182-C189, C199|LargeIntestine|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C180, C182-C189, C199|LargeIntestine|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C180, C182-C189, C199|LargeIntestine|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C180, C182-C189, C199|LargeIntestine|880|Sarcoma|8800/3|Sarcoma
C180, C182-C189, C199|LargeIntestine|880|Sarcoma|8801/3|SpindleCellSarcoma
C180, C182-C189, C199|LargeIntestine|880|Sarcoma|8802/3|GiantCellSarcoma
C180, C182-C189, C199|LargeIntestine|880|Sarcoma|8803/3|SmallCellSarcoma
C180, C182-C189, C199|LargeIntestine|880|Sarcoma|8804/3|SarcomaEpithelioid
C180, C182-C189, C199|LargeIntestine|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C180, C182-C189, C199|LargeIntestine|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C180, C182-C189, C199|LargeIntestine|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C180, C182-C189, C199|LargeIntestine|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C180, C182-C189, C199|LargeIntestine|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C180, C182-C189, C199|LargeIntestine|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C180, C182-C189, C199|LargeIntestine|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C180, C182-C189, C199|LargeIntestine|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C180, C182-C189, C199|LargeIntestine|885|Liposarcoma|8850/3|Liposarcoma
C180, C182-C189, C199|LargeIntestine|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C180, C182-C189, C199|LargeIntestine|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C180, C182-C189, C199|LargeIntestine|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C180, C182-C189, C199|LargeIntestine|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C180, C182-C189, C199|LargeIntestine|885|Liposarcoma|8855/3|Liposarcoma
C180, C182-C189, C199|LargeIntestine|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C180, C182-C189, C199|LargeIntestine|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C180, C182-C189, C199|LargeIntestine|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C180, C182-C189, C199|LargeIntestine|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C180, C182-C189, C199|LargeIntestine|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C180, C182-C189, C199|LargeIntestine|889|MyomatousNeoplasm|8895/3|Myosarcoma
C180, C182-C189, C199|LargeIntestine|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C180, C182-C189, C199|LargeIntestine|893|StromalSarcoma|8934/3|Carcinofibroma
C180, C182-C189, C199|LargeIntestine|893|StromalSarcoma|8935/3|StromalSarcoma
C180, C182-C189, C199|LargeIntestine|893|StromalSarcoma|8936/3|HighRiskGastrointestinalStromalTumor
C180, C182-C189, C199|LargeIntestine|898|Carcinosarcoma|8980/3|Carcinosarcoma
C180, C182-C189, C199|LargeIntestine|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C180, C182-C189, C199|LargeIntestine|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C180, C182-C189, C199|LargeIntestine|959|Lymphoma|9590/3|Lymphoma
C180, C182-C189, C199|LargeIntestine|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C180, C182-C189, C199|LargeIntestine|959|Lymphoma|9596/3|CompositeLymphoma
C180, C182-C189, C199|LargeIntestine|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C180, C182-C189, C199|LargeIntestine|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C180, C182-C189, C199|LargeIntestine|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C180, C182-C189, C199|LargeIntestine|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C180, C182-C189, C199|LargeIntestine|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C180, C182-C189, C199|LargeIntestine|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C180, C182-C189, C199|LargeIntestine|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C180, C182-C189, C199|LargeIntestine|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C180, C182-C189, C199|LargeIntestine|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C180, C182-C189, C199|LargeIntestine|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C180, C182-C189, C199|LargeIntestine|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C180, C182-C189, C199|LargeIntestine|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C180, C182-C189, C199|LargeIntestine|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C180, C182-C189, C199|LargeIntestine|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C180, C182-C189, C199|LargeIntestine|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C180, C182-C189, C199|LargeIntestine|967|BCellLymphomas|9673/3|MantleCellLymphoma
C180, C182-C189, C199|LargeIntestine|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C180, C182-C189, C199|LargeIntestine|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C180, C182-C189, C199|LargeIntestine|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C180, C182-C189, C199|LargeIntestine|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C180, C182-C189, C199|LargeIntestine|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C180, C182-C189, C199|LargeIntestine|969|FollicularAdenoma|9690/3|LymphomaFollicular
C180, C182-C189, C199|LargeIntestine|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C180, C182-C189, C199|LargeIntestine|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C180, C182-C189, C199|LargeIntestine|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C180, C182-C189, C199|LargeIntestine|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C180, C182-C189, C199|LargeIntestine|970|TCellLymphoma|9701/3|SezarySyndrome
C180, C182-C189, C199|LargeIntestine|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C180, C182-C189, C199|LargeIntestine|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C180, C182-C189, C199|LargeIntestine|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C180, C182-C189, C199|LargeIntestine|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C180, C182-C189, C199|LargeIntestine|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C180, C182-C189, C199|LargeIntestine|971|AdultNonHodgkinLymphoma|9717/3|IntestinalTCellLymphomaNOS
C180, C182-C189, C199|LargeIntestine|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C180, C182-C189, C199|LargeIntestine|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C180, C182-C189, C199|LargeIntestine|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C180, C182-C189, C199|LargeIntestine|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C180, C182-C189, C199|LargeIntestine|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C180, C182-C189, C199|LargeIntestine|973|Plasmacytoma|9731/3|Plasmacytoma
C180, C182-C189, C199|LargeIntestine|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C180, C182-C189, C199|LargeIntestine|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C180, C182-C189, C199|LargeIntestine|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C180, C182-C189, C199|LargeIntestine|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C180, C182-C189, C199|LargeIntestine|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C180, C182-C189, C199|LargeIntestine|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C180, C182-C189, C199|LargeIntestine|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C180, C182-C189, C199|LargeIntestine|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C180, C182-C189, C199|LargeIntestine|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C180, C182-C189, C199|LargeIntestine|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C180, C182-C189, C199|LargeIntestine|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C180, C182-C189, C199|LargeIntestine|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C180, C182-C189, C199|LargeIntestine|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C180, C182-C189, C199|LargeIntestine|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C180, C182-C189, C199|LargeIntestine|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C180, C182-C189, C199|LargeIntestine|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9812/3|null
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9813/3|null
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9814/3|null
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9817/3|null
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9818/3|null
C180, C182-C189, C199|LargeIntestine|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C180, C182-C189, C199|LargeIntestine|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C180, C182-C189, C199|LargeIntestine|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C180, C182-C189, C199|LargeIntestine|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C180, C182-C189, C199|LargeIntestine|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C180, C182-C189, C199|LargeIntestine|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C180, C182-C189, C199|LargeIntestine|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C180, C182-C189, C199|LargeIntestine|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C181|Appendix|801|Carcinoma|8010/2|InSituCancer
C181|Appendix|801|Carcinoma|8010/3|CarcinomaNOSDNE
C181|Appendix|801|Carcinoma|8011/3|MalignantEpithelioma
C181|Appendix|801|Carcinoma|8012/3|LargeCellCarcinoma
C181|Appendix|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C181|Appendix|801|Carcinoma|8014/3|LargeCellCarcinoma
C181|Appendix|801|Carcinoma|8015/3|GlassyCellCarcinoma
C181|Appendix|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C181|Appendix|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C181|Appendix|802|Carcinoma|8022/3|PleomorphicCarcinoma
C181|Appendix|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C181|Appendix|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C181|Appendix|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C181|Appendix|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C181|Appendix|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C181|Appendix|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C181|Appendix|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C181|Appendix|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C181|Appendix|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C181|Appendix|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C181|Appendix|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C181|Appendix|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C181|Appendix|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C181|Appendix|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C181|Appendix|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C181|Appendix|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C181|Appendix|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C181|Appendix|814|Adenocarcinoma|8140/3|Adenocarcinoma
C181|Appendix|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C181|Appendix|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C181|Appendix|814|Adenocarcinoma|8145/3|DiffuseTypeAdenocarcinoma
C181|Appendix|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C181|Appendix|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C181|Appendix|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C181|Appendix|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C181|Appendix|822|FamilialAdenomatousPolyposis|8220/2|AdenocarcinomaInSitu
C181|Appendix|822|FamilialAdenomatousPolyposis|8220/3|FamilialAdenomatousPolyposis
C181|Appendix|822|FamilialAdenomatousPolyposis|8221/2|AdenomatousPolyp
C181|Appendix|822|FamilialAdenomatousPolyposis|8221/3|AdenomatousPolyp
C181|Appendix|823|SolidCarcinoma|8230/2|InSituCancer
C181|Appendix|823|SolidCarcinoma|8230/3|SolidCarcinoma
C181|Appendix|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C181|Appendix|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C181|Appendix|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C181|Appendix|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C181|Appendix|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C181|Appendix|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C181|Appendix|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C181|Appendix|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C181|Appendix|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C181|Appendix|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C181|Appendix|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C181|Appendix|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C181|Appendix|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C181|Appendix|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C181|Appendix|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C181|Appendix|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C181|Appendix|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C181|Appendix|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C181|Appendix|847|MucinousCystadenocarcinoma|8470/2|MucinousCystadenocarcinoma
C181|Appendix|847|MucinousCystadenocarcinoma|8470/3|MucinousCystadenocarcinoma
C181|Appendix|847|MucinousCystadenocarcinoma|8471/3|PapillaryMucinousCystadenocarcinoma
C181|Appendix|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C181|Appendix|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C181|Appendix|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C181|Appendix|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C181|Appendix|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C181|Appendix|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C181|Appendix|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C181|Appendix|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C181|Appendix|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C181|Appendix|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C181|Appendix|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C181|Appendix|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C181|Appendix|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C181|Appendix|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C181|Appendix|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C181|Appendix|880|Sarcoma|8800/3|Sarcoma
C181|Appendix|880|Sarcoma|8801/3|SpindleCellSarcoma
C181|Appendix|880|Sarcoma|8802/3|GiantCellSarcoma
C181|Appendix|880|Sarcoma|8803/3|SmallCellSarcoma
C181|Appendix|880|Sarcoma|8804/3|SarcomaEpithelioid
C181|Appendix|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C181|Appendix|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C181|Appendix|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C181|Appendix|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C181|Appendix|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C181|Appendix|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C181|Appendix|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C181|Appendix|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C181|Appendix|885|Liposarcoma|8850/3|Liposarcoma
C181|Appendix|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C181|Appendix|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C181|Appendix|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C181|Appendix|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C181|Appendix|885|Liposarcoma|8855/3|Liposarcoma
C181|Appendix|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C181|Appendix|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C181|Appendix|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C181|Appendix|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C181|Appendix|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C181|Appendix|889|MyomatousNeoplasm|8895/3|Myosarcoma
C181|Appendix|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C181|Appendix|893|StromalSarcoma|8934/3|Carcinofibroma
C181|Appendix|893|StromalSarcoma|8935/3|StromalSarcoma
C181|Appendix|893|StromalSarcoma|8936/3|HighRiskGastrointestinalStromalTumor
C181|Appendix|898|Carcinosarcoma|8980/3|Carcinosarcoma
C181|Appendix|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C181|Appendix|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C181|Appendix|959|Lymphoma|9590/3|Lymphoma
C181|Appendix|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C181|Appendix|959|Lymphoma|9596/3|CompositeLymphoma
C181|Appendix|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C181|Appendix|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C181|Appendix|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C181|Appendix|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C181|Appendix|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C181|Appendix|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C181|Appendix|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C181|Appendix|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C181|Appendix|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C181|Appendix|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C181|Appendix|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C181|Appendix|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C181|Appendix|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C181|Appendix|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C181|Appendix|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C181|Appendix|967|BCellLymphomas|9673/3|MantleCellLymphoma
C181|Appendix|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C181|Appendix|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C181|Appendix|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C181|Appendix|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C181|Appendix|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C181|Appendix|969|FollicularAdenoma|9690/3|LymphomaFollicular
C181|Appendix|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C181|Appendix|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C181|Appendix|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C181|Appendix|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C181|Appendix|970|TCellLymphoma|9701/3|SezarySyndrome
C181|Appendix|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C181|Appendix|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C181|Appendix|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C181|Appendix|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C181|Appendix|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C181|Appendix|971|AdultNonHodgkinLymphoma|9717/3|IntestinalTCellLymphomaNOS
C181|Appendix|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C181|Appendix|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C181|Appendix|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C181|Appendix|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C181|Appendix|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C181|Appendix|973|Plasmacytoma|9731/3|Plasmacytoma
C181|Appendix|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C181|Appendix|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C181|Appendix|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C181|Appendix|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C181|Appendix|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C181|Appendix|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C181|Appendix|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C181|Appendix|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C181|Appendix|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C181|Appendix|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C181|Appendix|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C181|Appendix|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C181|Appendix|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C181|Appendix|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C181|Appendix|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C181|Appendix|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C181|Appendix|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C181|Appendix|981|PrecursorLymphoidNeoplasm|9812/3|null
C181|Appendix|981|PrecursorLymphoidNeoplasm|9813/3|null
C181|Appendix|981|PrecursorLymphoidNeoplasm|9814/3|null
C181|Appendix|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C181|Appendix|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C181|Appendix|981|PrecursorLymphoidNeoplasm|9817/3|null
C181|Appendix|981|PrecursorLymphoidNeoplasm|9818/3|null
C181|Appendix|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C181|Appendix|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C181|Appendix|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C181|Appendix|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C181|Appendix|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C181|Appendix|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C181|Appendix|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C181|Appendix|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C209|Rectal|801|Carcinoma|8010/2|InSituCancer
C209|Rectal|801|Carcinoma|8010/3|CarcinomaNOSDNE
C209|Rectal|801|Carcinoma|8011/3|MalignantEpithelioma
C209|Rectal|801|Carcinoma|8012/3|LargeCellCarcinoma
C209|Rectal|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C209|Rectal|801|Carcinoma|8014/3|LargeCellCarcinoma
C209|Rectal|801|Carcinoma|8015/3|GlassyCellCarcinoma
C209|Rectal|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C209|Rectal|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C209|Rectal|802|Carcinoma|8022/3|PleomorphicCarcinoma
C209|Rectal|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C209|Rectal|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C209|Rectal|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C209|Rectal|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C209|Rectal|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C209|Rectal|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C209|Rectal|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C209|Rectal|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C209|Rectal|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C209|Rectal|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C209|Rectal|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C209|Rectal|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C209|Rectal|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C209|Rectal|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C209|Rectal|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C209|Rectal|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C209|Rectal|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C209|Rectal|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C209|Rectal|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C209|Rectal|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C209|Rectal|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C209|Rectal|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C209|Rectal|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C209|Rectal|814|Adenocarcinoma|8140/3|Adenocarcinoma
C209|Rectal|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C209|Rectal|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C209|Rectal|814|Adenocarcinoma|8145/3|DiffuseTypeAdenocarcinoma
C209|Rectal|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C209|Rectal|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C209|Rectal|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C209|Rectal|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C209|Rectal|821|AdenocarcinomaInAdenomatousPolyp|8213/3|SerratedAdenocarcinoma
C209|Rectal|822|FamilialAdenomatousPolyposis|8220/2|AdenocarcinomaInSitu
C209|Rectal|822|FamilialAdenomatousPolyposis|8220/3|FamilialAdenomatousPolyposis
C209|Rectal|822|FamilialAdenomatousPolyposis|8221/2|AdenomatousPolyp
C209|Rectal|822|FamilialAdenomatousPolyposis|8221/3|AdenomatousPolyp
C209|Rectal|823|SolidCarcinoma|8230/2|InSituCancer
C209|Rectal|823|SolidCarcinoma|8230/3|SolidCarcinoma
C209|Rectal|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C209|Rectal|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C209|Rectal|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C209|Rectal|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C209|Rectal|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C209|Rectal|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C209|Rectal|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C209|Rectal|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C209|Rectal|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C209|Rectal|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C209|Rectal|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C209|Rectal|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C209|Rectal|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C209|Rectal|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C209|Rectal|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C209|Rectal|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C209|Rectal|826|PapillaryAdenocarcinoma|8265/3|MicropapillaryCarcinoma
C209|Rectal|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C209|Rectal|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C209|Rectal|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C209|Rectal|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C209|Rectal|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C209|Rectal|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C209|Rectal|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C209|Rectal|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C209|Rectal|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C209|Rectal|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C209|Rectal|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C209|Rectal|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C209|Rectal|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C209|Rectal|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C209|Rectal|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C209|Rectal|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C209|Rectal|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C209|Rectal|872|Melanoma|8720/2|Stage0SkinMelanoma
C209|Rectal|872|Melanoma|8720/3|Melanoma
C209|Rectal|872|Melanoma|8721/3|NodularMelanoma
C209|Rectal|872|Melanoma|8722/3|BalloonCellMelanoma
C209|Rectal|872|Melanoma|8723/3|RegressingMelanoma
C209|Rectal|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C209|Rectal|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C209|Rectal|874|Nevus|8745/3|DesmoplasticMelanoma
C209|Rectal|874|Nevus|8746/3|MucosalLentiginousMelanoma
C209|Rectal|876|Nevus|8761/3|GiantCongenitalNevus
C209|Rectal|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C209|Rectal|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C209|Rectal|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C209|Rectal|880|Sarcoma|8800/3|Sarcoma
C209|Rectal|880|Sarcoma|8801/3|SpindleCellSarcoma
C209|Rectal|880|Sarcoma|8802/3|GiantCellSarcoma
C209|Rectal|880|Sarcoma|8803/3|SmallCellSarcoma
C209|Rectal|880|Sarcoma|8804/3|SarcomaEpithelioid
C209|Rectal|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C209|Rectal|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C209|Rectal|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C209|Rectal|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C209|Rectal|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C209|Rectal|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C209|Rectal|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C209|Rectal|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C209|Rectal|885|Liposarcoma|8850/3|Liposarcoma
C209|Rectal|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C209|Rectal|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C209|Rectal|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C209|Rectal|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C209|Rectal|885|Liposarcoma|8855/3|Liposarcoma
C209|Rectal|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C209|Rectal|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C209|Rectal|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C209|Rectal|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C209|Rectal|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C209|Rectal|889|MyomatousNeoplasm|8895/3|Myosarcoma
C209|Rectal|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C209|Rectal|893|StromalSarcoma|8934/3|Carcinofibroma
C209|Rectal|893|StromalSarcoma|8935/3|StromalSarcoma
C209|Rectal|893|StromalSarcoma|8936/3|HighRiskGastrointestinalStromalTumor
C209|Rectal|898|Carcinosarcoma|8980/3|Carcinosarcoma
C209|Rectal|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C209|Rectal|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C209|Rectal|959|Lymphoma|9590/3|Lymphoma
C209|Rectal|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C209|Rectal|959|Lymphoma|9596/3|CompositeLymphoma
C209|Rectal|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C209|Rectal|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C209|Rectal|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C209|Rectal|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C209|Rectal|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C209|Rectal|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C209|Rectal|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C209|Rectal|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C209|Rectal|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C209|Rectal|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C209|Rectal|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C209|Rectal|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C209|Rectal|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C209|Rectal|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C209|Rectal|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C209|Rectal|967|BCellLymphomas|9673/3|MantleCellLymphoma
C209|Rectal|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C209|Rectal|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C209|Rectal|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C209|Rectal|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C209|Rectal|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C209|Rectal|969|FollicularAdenoma|9690/3|LymphomaFollicular
C209|Rectal|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C209|Rectal|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C209|Rectal|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C209|Rectal|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C209|Rectal|970|TCellLymphoma|9701/3|SezarySyndrome
C209|Rectal|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C209|Rectal|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C209|Rectal|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C209|Rectal|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C209|Rectal|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C209|Rectal|971|AdultNonHodgkinLymphoma|9717/3|IntestinalTCellLymphomaNOS
C209|Rectal|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C209|Rectal|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C209|Rectal|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C209|Rectal|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C209|Rectal|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C209|Rectal|973|Plasmacytoma|9731/3|Plasmacytoma
C209|Rectal|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C209|Rectal|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C209|Rectal|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C209|Rectal|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C209|Rectal|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C209|Rectal|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C209|Rectal|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C209|Rectal|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C209|Rectal|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C209|Rectal|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C209|Rectal|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C209|Rectal|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C209|Rectal|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C209|Rectal|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C209|Rectal|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C209|Rectal|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C209|Rectal|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C209|Rectal|981|PrecursorLymphoidNeoplasm|9812/3|null
C209|Rectal|981|PrecursorLymphoidNeoplasm|9813/3|null
C209|Rectal|981|PrecursorLymphoidNeoplasm|9814/3|null
C209|Rectal|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C209|Rectal|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C209|Rectal|981|PrecursorLymphoidNeoplasm|9817/3|null
C209|Rectal|981|PrecursorLymphoidNeoplasm|9818/3|null
C209|Rectal|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C209|Rectal|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C209|Rectal|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C209|Rectal|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C209|Rectal|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C209|Rectal|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C209|Rectal|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C209|Rectal|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C210-C212,C218|AnalCanal|801|Carcinoma|8010/2|InSituCancer
C210-C212,C218|AnalCanal|801|Carcinoma|8010/3|CarcinomaNOSDNE
C210-C212,C218|AnalCanal|801|Carcinoma|8011/3|MalignantEpithelioma
C210-C212,C218|AnalCanal|801|Carcinoma|8012/3|LargeCellCarcinoma
C210-C212,C218|AnalCanal|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C210-C212,C218|AnalCanal|801|Carcinoma|8014/3|LargeCellCarcinoma
C210-C212,C218|AnalCanal|801|Carcinoma|8015/3|GlassyCellCarcinoma
C210-C212,C218|AnalCanal|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C210-C212,C218|AnalCanal|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C210-C212,C218|AnalCanal|802|Carcinoma|8022/3|PleomorphicCarcinoma
C210-C212,C218|AnalCanal|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C210-C212,C218|AnalCanal|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C210-C212,C218|AnalCanal|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C210-C212,C218|AnalCanal|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C210-C212,C218|AnalCanal|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C210-C212,C218|AnalCanal|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C210-C212,C218|AnalCanal|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C210-C212,C218|AnalCanal|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8077/2|IntraepithelialNeoplasia
C210-C212,C218|AnalCanal|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C210-C212,C218|AnalCanal|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C210-C212,C218|AnalCanal|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C210-C212,C218|AnalCanal|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C210-C212,C218|AnalCanal|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C210-C212,C218|AnalCanal|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C210-C212,C218|AnalCanal|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C210-C212,C218|AnalCanal|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C210-C212,C218|AnalCanal|814|Adenocarcinoma|8140/3|Adenocarcinoma
C210-C212,C218|AnalCanal|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C210-C212,C218|AnalCanal|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C210-C212,C218|AnalCanal|814|Adenocarcinoma|8145/3|DiffuseTypeAdenocarcinoma
C210-C212,C218|AnalCanal|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C210-C212,C218|AnalCanal|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C210-C212,C218|AnalCanal|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C210-C212,C218|AnalCanal|821|AdenocarcinomaInAdenomatousPolyp|8215/3|AnalGlandsAdenocarcinoma
C210-C212,C218|AnalCanal|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C210-C212,C218|AnalCanal|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C210-C212,C218|AnalCanal|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C210-C212,C218|AnalCanal|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C210-C212,C218|AnalCanal|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C210-C212,C218|AnalCanal|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C210-C212,C218|AnalCanal|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C210-C212,C218|AnalCanal|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C210-C212,C218|AnalCanal|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C210-C212,C218|AnalCanal|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C210-C212,C218|AnalCanal|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C210-C212,C218|AnalCanal|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C210-C212,C218|AnalCanal|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C210-C212,C218|AnalCanal|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C210-C212,C218|AnalCanal|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C210-C212,C218|AnalCanal|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C210-C212,C218|AnalCanal|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C210-C212,C218|AnalCanal|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C210-C212,C218|AnalCanal|850|DuctalCarcinoma|8500/2|DuctalBreastCarcinomaInSitu
C210-C212,C218|AnalCanal|850|DuctalCarcinoma|8500/3|InvasiveBreastCarcinoma
C210-C212,C218|AnalCanal|850|DuctalCarcinoma|8503/2|IntraductalPapillaryBreastCarcinoma
C210-C212,C218|AnalCanal|850|DuctalCarcinoma|8503/3|IntraductalPapillaryBreastCarcinoma
C210-C212,C218|AnalCanal|850|DuctalCarcinoma|8504/2|IntracysticPapillaryBreastCarcinoma
C210-C212,C218|AnalCanal|850|DuctalCarcinoma|8504/3|IntracysticPapillaryBreastCarcinoma
C210-C212,C218|AnalCanal|854|PagetDiseaseExtramammary|8542/3|PagetDiseaseExtramammary
C210-C212,C218|AnalCanal|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C210-C212,C218|AnalCanal|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C210-C212,C218|AnalCanal|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C210-C212,C218|AnalCanal|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C210-C212,C218|AnalCanal|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C210-C212,C218|AnalCanal|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C210-C212,C218|AnalCanal|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C210-C212,C218|AnalCanal|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C210-C212,C218|AnalCanal|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C210-C212,C218|AnalCanal|872|Melanoma|8720/2|Stage0SkinMelanoma
C210-C212,C218|AnalCanal|872|Melanoma|8720/3|Melanoma
C210-C212,C218|AnalCanal|872|Melanoma|8721/3|NodularMelanoma
C210-C212,C218|AnalCanal|872|Melanoma|8722/3|BalloonCellMelanoma
C210-C212,C218|AnalCanal|872|Melanoma|8723/3|RegressingMelanoma
C210-C212,C218|AnalCanal|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C210-C212,C218|AnalCanal|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C210-C212,C218|AnalCanal|874|Nevus|8745/3|DesmoplasticMelanoma
C210-C212,C218|AnalCanal|874|Nevus|8746/3|MucosalLentiginousMelanoma
C210-C212,C218|AnalCanal|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C210-C212,C218|AnalCanal|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C210-C212,C218|AnalCanal|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C210-C212,C218|AnalCanal|880|Sarcoma|8800/3|Sarcoma
C210-C212,C218|AnalCanal|880|Sarcoma|8801/3|SpindleCellSarcoma
C210-C212,C218|AnalCanal|880|Sarcoma|8802/3|GiantCellSarcoma
C210-C212,C218|AnalCanal|880|Sarcoma|8803/3|SmallCellSarcoma
C210-C212,C218|AnalCanal|880|Sarcoma|8804/3|SarcomaEpithelioid
C210-C212,C218|AnalCanal|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C210-C212,C218|AnalCanal|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C210-C212,C218|AnalCanal|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C210-C212,C218|AnalCanal|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C210-C212,C218|AnalCanal|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C210-C212,C218|AnalCanal|889|MyomatousNeoplasm|8895/3|Myosarcoma
C210-C212,C218|AnalCanal|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C210-C212,C218|AnalCanal|959|Lymphoma|9590/3|Lymphoma
C210-C212,C218|AnalCanal|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C210-C212,C218|AnalCanal|959|Lymphoma|9596/3|CompositeLymphoma
C210-C212,C218|AnalCanal|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C210-C212,C218|AnalCanal|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C210-C212,C218|AnalCanal|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C210-C212,C218|AnalCanal|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C210-C212,C218|AnalCanal|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C210-C212,C218|AnalCanal|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C210-C212,C218|AnalCanal|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C210-C212,C218|AnalCanal|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C210-C212,C218|AnalCanal|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C210-C212,C218|AnalCanal|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C210-C212,C218|AnalCanal|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C210-C212,C218|AnalCanal|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C210-C212,C218|AnalCanal|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C210-C212,C218|AnalCanal|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C210-C212,C218|AnalCanal|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C210-C212,C218|AnalCanal|967|BCellLymphomas|9673/3|MantleCellLymphoma
C210-C212,C218|AnalCanal|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C210-C212,C218|AnalCanal|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C210-C212,C218|AnalCanal|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C210-C212,C218|AnalCanal|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C210-C212,C218|AnalCanal|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C210-C212,C218|AnalCanal|969|FollicularAdenoma|9690/3|LymphomaFollicular
C210-C212,C218|AnalCanal|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C210-C212,C218|AnalCanal|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C210-C212,C218|AnalCanal|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C210-C212,C218|AnalCanal|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C210-C212,C218|AnalCanal|970|TCellLymphoma|9701/3|SezarySyndrome
C210-C212,C218|AnalCanal|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C210-C212,C218|AnalCanal|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C210-C212,C218|AnalCanal|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C210-C212,C218|AnalCanal|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C210-C212,C218|AnalCanal|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C210-C212,C218|AnalCanal|971|AdultNonHodgkinLymphoma|9717/3|IntestinalTCellLymphomaNOS
C210-C212,C218|AnalCanal|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C210-C212,C218|AnalCanal|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C210-C212,C218|AnalCanal|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C210-C212,C218|AnalCanal|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C210-C212,C218|AnalCanal|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C210-C212,C218|AnalCanal|973|Plasmacytoma|9731/3|Plasmacytoma
C210-C212,C218|AnalCanal|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C210-C212,C218|AnalCanal|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C210-C212,C218|AnalCanal|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C210-C212,C218|AnalCanal|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C210-C212,C218|AnalCanal|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C210-C212,C218|AnalCanal|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C210-C212,C218|AnalCanal|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C210-C212,C218|AnalCanal|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C210-C212,C218|AnalCanal|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C210-C212,C218|AnalCanal|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C210-C212,C218|AnalCanal|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C210-C212,C218|AnalCanal|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C210-C212,C218|AnalCanal|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C210-C212,C218|AnalCanal|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C210-C212,C218|AnalCanal|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C210-C212,C218|AnalCanal|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9812/3|null
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9813/3|null
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9814/3|null
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9817/3|null
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9818/3|null
C210-C212,C218|AnalCanal|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C210-C212,C218|AnalCanal|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C210-C212,C218|AnalCanal|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C210-C212,C218|AnalCanal|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C210-C212,C218|AnalCanal|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C210-C212,C218|AnalCanal|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C210-C212,C218|AnalCanal|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C210-C212,C218|AnalCanal|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C220|Liver|801|Carcinoma|8010/2|InSituCancer
C220|Liver|801|Carcinoma|8010/3|CarcinomaNOSDNE
C220|Liver|801|Carcinoma|8011/3|MalignantEpithelioma
C220|Liver|801|Carcinoma|8012/3|LargeCellCarcinoma
C220|Liver|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C220|Liver|801|Carcinoma|8014/3|LargeCellCarcinoma
C220|Liver|801|Carcinoma|8015/3|GlassyCellCarcinoma
C220|Liver|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C220|Liver|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C220|Liver|802|Carcinoma|8022/3|PleomorphicCarcinoma
C220|Liver|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C220|Liver|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C220|Liver|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C220|Liver|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C220|Liver|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C220|Liver|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C220|Liver|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C220|Liver|814|Adenocarcinoma|8140/3|Adenocarcinoma
C220|Liver|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C220|Liver|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C220|Liver|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C220|Liver|816|Cholangiocarcinoma|8160/3|Cholangiocarcinoma
C220|Liver|816|Cholangiocarcinoma|8161/3|BileDuctCystadenocarcinoma
C220|Liver|817|HepatocellularCarcinoma|8170/3|HepatocellularCarcinoma
C220|Liver|817|HepatocellularCarcinoma|8171/3|FibrolamellarCarcinoma
C220|Liver|817|HepatocellularCarcinoma|8172/3|ScirrhousHepatocellularCarcinoma
C220|Liver|817|HepatocellularCarcinoma|8173/3|HepatocellularCarcinoma
C220|Liver|817|HepatocellularCarcinoma|8174/3|HepatocellularCarcinoma
C220|Liver|817|HepatocellularCarcinoma|8175/3|HepatocellularCarcinoma
C220|Liver|818|IntrahepaticCholangiocarcinoma|8180/3|Cholangiocarcinoma
C220|Liver|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C220|Liver|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C220|Liver|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C220|Liver|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C220|Liver|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C220|Liver|850|DuctalCarcinoma|8500/2|DuctalBreastCarcinomaInSitu
C220|Liver|850|DuctalCarcinoma|8500/3|InvasiveBreastCarcinoma
C220|Liver|850|DuctalCarcinoma|8501/2|Comedocarcinoma
C220|Liver|850|DuctalCarcinoma|8501/3|Comedocarcinoma
C220|Liver|850|DuctalCarcinoma|8503/2|IntraductalPapillaryBreastCarcinoma
C220|Liver|850|DuctalCarcinoma|8503/3|IntraductalPapillaryBreastCarcinoma
C220|Liver|850|DuctalCarcinoma|8504/2|IntracysticPapillaryBreastCarcinoma
C220|Liver|850|DuctalCarcinoma|8504/3|IntracysticPapillaryBreastCarcinoma
C220|Liver|850|DuctalCarcinoma|8507/2|MicropapillaryCarcinoma
C220|Liver|850|DuctalCarcinoma|8508/3|SecretoryBreastCarcinoma
C220|Liver|880|Sarcoma|8800/3|Sarcoma
C220|Liver|880|Sarcoma|8801/3|SpindleCellSarcoma
C220|Liver|880|Sarcoma|8802/3|GiantCellSarcoma
C220|Liver|880|Sarcoma|8803/3|SmallCellSarcoma
C220|Liver|880|Sarcoma|8804/3|SarcomaEpithelioid
C220|Liver|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C220|Liver|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C220|Liver|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C220|Liver|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C220|Liver|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C220|Liver|889|MyomatousNeoplasm|8895/3|Myosarcoma
C220|Liver|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C220|Liver|897|Hepatoblastoma|8970/3|Hepatoblastoma
C220|Liver|898|Carcinosarcoma|8980/3|Carcinosarcoma
C220|Liver|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C220|Liver|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C220|Liver|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C220|Liver|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C220|Liver|912|NeoplasmsVascularTissue|9124/3|KupfferCellSarcoma
C220|Liver|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C220|Liver|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C220|Liver|959|Lymphoma|9590/3|Lymphoma
C220|Liver|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C220|Liver|959|Lymphoma|9596/3|CompositeLymphoma
C220|Liver|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C220|Liver|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C220|Liver|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C220|Liver|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C220|Liver|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C220|Liver|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C220|Liver|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C220|Liver|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C220|Liver|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C220|Liver|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C220|Liver|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C220|Liver|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C220|Liver|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C220|Liver|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C220|Liver|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C220|Liver|967|BCellLymphomas|9673/3|MantleCellLymphoma
C220|Liver|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C220|Liver|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C220|Liver|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C220|Liver|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C220|Liver|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C220|Liver|969|FollicularAdenoma|9690/3|LymphomaFollicular
C220|Liver|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C220|Liver|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C220|Liver|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C220|Liver|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C220|Liver|970|TCellLymphoma|9701/3|SezarySyndrome
C220|Liver|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C220|Liver|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C220|Liver|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C220|Liver|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C220|Liver|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C220|Liver|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C220|Liver|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C220|Liver|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C220|Liver|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C220|Liver|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C220|Liver|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C220|Liver|973|Plasmacytoma|9731/3|Plasmacytoma
C220|Liver|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C220|Liver|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C220|Liver|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C220|Liver|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C220|Liver|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C220|Liver|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C220|Liver|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C220|Liver|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C220|Liver|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C220|Liver|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C220|Liver|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C220|Liver|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C220|Liver|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C220|Liver|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C220|Liver|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C220|Liver|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C220|Liver|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C220|Liver|981|PrecursorLymphoidNeoplasm|9812/3|null
C220|Liver|981|PrecursorLymphoidNeoplasm|9813/3|null
C220|Liver|981|PrecursorLymphoidNeoplasm|9814/3|null
C220|Liver|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C220|Liver|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C220|Liver|981|PrecursorLymphoidNeoplasm|9817/3|null
C220|Liver|981|PrecursorLymphoidNeoplasm|9818/3|null
C220|Liver|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C220|Liver|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C220|Liver|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C220|Liver|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C220|Liver|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C220|Liver|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C220|Liver|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C220|Liver|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C221|IntrahepaticBileDuct|801|Carcinoma|8010/2|InSituCancer
C221|IntrahepaticBileDuct|801|Carcinoma|8010/3|CarcinomaNOSDNE
C221|IntrahepaticBileDuct|801|Carcinoma|8011/3|MalignantEpithelioma
C221|IntrahepaticBileDuct|801|Carcinoma|8012/3|LargeCellCarcinoma
C221|IntrahepaticBileDuct|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C221|IntrahepaticBileDuct|801|Carcinoma|8014/3|LargeCellCarcinoma
C221|IntrahepaticBileDuct|801|Carcinoma|8015/3|GlassyCellCarcinoma
C221|IntrahepaticBileDuct|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C221|IntrahepaticBileDuct|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C221|IntrahepaticBileDuct|802|Carcinoma|8022/3|PleomorphicCarcinoma
C221|IntrahepaticBileDuct|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C221|IntrahepaticBileDuct|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C221|IntrahepaticBileDuct|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C221|IntrahepaticBileDuct|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C221|IntrahepaticBileDuct|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C221|IntrahepaticBileDuct|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C221|IntrahepaticBileDuct|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C221|IntrahepaticBileDuct|814|Adenocarcinoma|8140/3|Adenocarcinoma
C221|IntrahepaticBileDuct|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C221|IntrahepaticBileDuct|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C221|IntrahepaticBileDuct|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C221|IntrahepaticBileDuct|816|Cholangiocarcinoma|8160/3|Cholangiocarcinoma
C221|IntrahepaticBileDuct|816|Cholangiocarcinoma|8161/3|BileDuctCystadenocarcinoma
C221|IntrahepaticBileDuct|816|Cholangiocarcinoma|8162/3|HilarCholangiocarcinoma
C221|IntrahepaticBileDuct|817|HepatocellularCarcinoma|8170/3|HepatocellularCarcinoma
C221|IntrahepaticBileDuct|817|HepatocellularCarcinoma|8171/3|FibrolamellarCarcinoma
C221|IntrahepaticBileDuct|817|HepatocellularCarcinoma|8172/3|ScirrhousHepatocellularCarcinoma
C221|IntrahepaticBileDuct|817|HepatocellularCarcinoma|8173/3|HepatocellularCarcinoma
C221|IntrahepaticBileDuct|817|HepatocellularCarcinoma|8174/3|HepatocellularCarcinoma
C221|IntrahepaticBileDuct|817|HepatocellularCarcinoma|8175/3|HepatocellularCarcinoma
C221|IntrahepaticBileDuct|818|IntrahepaticCholangiocarcinoma|8180/3|Cholangiocarcinoma
C221|IntrahepaticBileDuct|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C221|IntrahepaticBileDuct|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C221|IntrahepaticBileDuct|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C221|IntrahepaticBileDuct|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C221|IntrahepaticBileDuct|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8500/2|DuctalBreastCarcinomaInSitu
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8500/3|InvasiveBreastCarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8501/2|Comedocarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8501/3|Comedocarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8503/2|IntraductalPapillaryBreastCarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8503/3|IntraductalPapillaryBreastCarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8504/2|IntracysticPapillaryBreastCarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8504/3|IntracysticPapillaryBreastCarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8507/2|MicropapillaryCarcinoma
C221|IntrahepaticBileDuct|850|DuctalCarcinoma|8508/3|SecretoryBreastCarcinoma
C221|IntrahepaticBileDuct|880|Sarcoma|8800/3|Sarcoma
C221|IntrahepaticBileDuct|880|Sarcoma|8801/3|SpindleCellSarcoma
C221|IntrahepaticBileDuct|880|Sarcoma|8802/3|GiantCellSarcoma
C221|IntrahepaticBileDuct|880|Sarcoma|8803/3|SmallCellSarcoma
C221|IntrahepaticBileDuct|880|Sarcoma|8804/3|SarcomaEpithelioid
C221|IntrahepaticBileDuct|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C221|IntrahepaticBileDuct|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C221|IntrahepaticBileDuct|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C221|IntrahepaticBileDuct|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C221|IntrahepaticBileDuct|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C221|IntrahepaticBileDuct|889|MyomatousNeoplasm|8895/3|Myosarcoma
C221|IntrahepaticBileDuct|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C221|IntrahepaticBileDuct|898|Carcinosarcoma|8980/3|Carcinosarcoma
C221|IntrahepaticBileDuct|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C221|IntrahepaticBileDuct|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C221|IntrahepaticBileDuct|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C221|IntrahepaticBileDuct|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C221|IntrahepaticBileDuct|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C221|IntrahepaticBileDuct|959|Lymphoma|9590/3|Lymphoma
C221|IntrahepaticBileDuct|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C221|IntrahepaticBileDuct|959|Lymphoma|9596/3|CompositeLymphoma
C221|IntrahepaticBileDuct|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C221|IntrahepaticBileDuct|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C221|IntrahepaticBileDuct|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C221|IntrahepaticBileDuct|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C221|IntrahepaticBileDuct|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C221|IntrahepaticBileDuct|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C221|IntrahepaticBileDuct|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C221|IntrahepaticBileDuct|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C221|IntrahepaticBileDuct|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C221|IntrahepaticBileDuct|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C221|IntrahepaticBileDuct|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C221|IntrahepaticBileDuct|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C221|IntrahepaticBileDuct|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C221|IntrahepaticBileDuct|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C221|IntrahepaticBileDuct|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C221|IntrahepaticBileDuct|967|BCellLymphomas|9673/3|MantleCellLymphoma
C221|IntrahepaticBileDuct|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C221|IntrahepaticBileDuct|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C221|IntrahepaticBileDuct|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C221|IntrahepaticBileDuct|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C221|IntrahepaticBileDuct|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C221|IntrahepaticBileDuct|969|FollicularAdenoma|9690/3|LymphomaFollicular
C221|IntrahepaticBileDuct|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C221|IntrahepaticBileDuct|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C221|IntrahepaticBileDuct|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C221|IntrahepaticBileDuct|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C221|IntrahepaticBileDuct|970|TCellLymphoma|9701/3|SezarySyndrome
C221|IntrahepaticBileDuct|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C221|IntrahepaticBileDuct|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C221|IntrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C221|IntrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C221|IntrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C221|IntrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C221|IntrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C221|IntrahepaticBileDuct|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C221|IntrahepaticBileDuct|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C221|IntrahepaticBileDuct|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C221|IntrahepaticBileDuct|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C221|IntrahepaticBileDuct|973|Plasmacytoma|9731/3|Plasmacytoma
C221|IntrahepaticBileDuct|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C221|IntrahepaticBileDuct|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C221|IntrahepaticBileDuct|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C221|IntrahepaticBileDuct|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C221|IntrahepaticBileDuct|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C221|IntrahepaticBileDuct|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C221|IntrahepaticBileDuct|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C221|IntrahepaticBileDuct|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C221|IntrahepaticBileDuct|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C221|IntrahepaticBileDuct|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C221|IntrahepaticBileDuct|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C221|IntrahepaticBileDuct|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C221|IntrahepaticBileDuct|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C221|IntrahepaticBileDuct|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C221|IntrahepaticBileDuct|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C221|IntrahepaticBileDuct|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9812/3|null
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9813/3|null
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9814/3|null
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9817/3|null
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9818/3|null
C221|IntrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C221|IntrahepaticBileDuct|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C221|IntrahepaticBileDuct|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C221|IntrahepaticBileDuct|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C221|IntrahepaticBileDuct|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C221|IntrahepaticBileDuct|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C221|IntrahepaticBileDuct|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C221|IntrahepaticBileDuct|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C239-C241,C248-C249|ExtrahepaticBileDuct|801|Carcinoma|8010/2|InSituCancer
C239-C241,C248-C249|ExtrahepaticBileDuct|801|Carcinoma|8010/3|CarcinomaNOSDNE
C239-C241,C248-C249|ExtrahepaticBileDuct|801|Carcinoma|8011/3|MalignantEpithelioma
C239-C241,C248-C249|ExtrahepaticBileDuct|801|Carcinoma|8012/3|LargeCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|801|Carcinoma|8014/3|LargeCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|801|Carcinoma|8015/3|GlassyCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C239-C241,C248-C249|ExtrahepaticBileDuct|802|Carcinoma|8022/3|PleomorphicCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C239-C241,C248-C249|ExtrahepaticBileDuct|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C239-C241,C248-C249|ExtrahepaticBileDuct|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C239-C241,C248-C249|ExtrahepaticBileDuct|814|Adenocarcinoma|8140/3|Adenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C239-C241,C248-C249|ExtrahepaticBileDuct|816|Cholangiocarcinoma|8160/3|Cholangiocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|816|Cholangiocarcinoma|8161/3|BileDuctCystadenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|816|Cholangiocarcinoma|8162/3|HilarCholangiocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|816|Cholangiocarcinoma|8163/3|PancreatobiliarytypeCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C239-C241,C248-C249|ExtrahepaticBileDuct|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C239-C241,C248-C249|ExtrahepaticBileDuct|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C239-C241,C248-C249|ExtrahepaticBileDuct|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C239-C241,C248-C249|ExtrahepaticBileDuct|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C239-C241,C248-C249|ExtrahepaticBileDuct|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8500/2|DuctalBreastCarcinomaInSitu
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8500/3|InvasiveBreastCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8501/2|Comedocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8501/3|Comedocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8503/2|IntraductalPapillaryBreastCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8503/3|IntraductalPapillaryBreastCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8504/2|IntracysticPapillaryBreastCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8504/3|IntracysticPapillaryBreastCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8507/2|MicropapillaryCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|850|DuctalCarcinoma|8508/3|SecretoryBreastCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C239-C241,C248-C249|ExtrahepaticBileDuct|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C239-C241,C248-C249|ExtrahepaticBileDuct|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C239-C241,C248-C249|ExtrahepaticBileDuct|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C239-C241,C248-C249|ExtrahepaticBileDuct|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C239-C241,C248-C249|ExtrahepaticBileDuct|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C239-C241,C248-C249|ExtrahepaticBileDuct|880|Sarcoma|8800/3|Sarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|880|Sarcoma|8801/3|SpindleCellSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|880|Sarcoma|8802/3|GiantCellSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|880|Sarcoma|8803/3|SmallCellSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|880|Sarcoma|8804/3|SarcomaEpithelioid
C239-C241,C248-C249|ExtrahepaticBileDuct|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C239-C241,C248-C249|ExtrahepaticBileDuct|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|889|MyomatousNeoplasm|8895/3|Myosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|898|Carcinosarcoma|8980/3|Carcinosarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C239-C241,C248-C249|ExtrahepaticBileDuct|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C239-C241,C248-C249|ExtrahepaticBileDuct|959|Lymphoma|9590/3|Lymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|959|Lymphoma|9596/3|CompositeLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C239-C241,C248-C249|ExtrahepaticBileDuct|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C239-C241,C248-C249|ExtrahepaticBileDuct|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C239-C241,C248-C249|ExtrahepaticBileDuct|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C239-C241,C248-C249|ExtrahepaticBileDuct|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C239-C241,C248-C249|ExtrahepaticBileDuct|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C239-C241,C248-C249|ExtrahepaticBileDuct|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C239-C241,C248-C249|ExtrahepaticBileDuct|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C239-C241,C248-C249|ExtrahepaticBileDuct|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C239-C241,C248-C249|ExtrahepaticBileDuct|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C239-C241,C248-C249|ExtrahepaticBileDuct|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|967|BCellLymphomas|9673/3|MantleCellLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|969|FollicularAdenoma|9690/3|LymphomaFollicular
C239-C241,C248-C249|ExtrahepaticBileDuct|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C239-C241,C248-C249|ExtrahepaticBileDuct|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C239-C241,C248-C249|ExtrahepaticBileDuct|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|970|TCellLymphoma|9701/3|SezarySyndrome
C239-C241,C248-C249|ExtrahepaticBileDuct|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C239-C241,C248-C249|ExtrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C239-C241,C248-C249|ExtrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C239-C241,C248-C249|ExtrahepaticBileDuct|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C239-C241,C248-C249|ExtrahepaticBileDuct|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C239-C241,C248-C249|ExtrahepaticBileDuct|973|Plasmacytoma|9731/3|Plasmacytoma
C239-C241,C248-C249|ExtrahepaticBileDuct|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C239-C241,C248-C249|ExtrahepaticBileDuct|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C239-C241,C248-C249|ExtrahepaticBileDuct|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C239-C241,C248-C249|ExtrahepaticBileDuct|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C239-C241,C248-C249|ExtrahepaticBileDuct|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C239-C241,C248-C249|ExtrahepaticBileDuct|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C239-C241,C248-C249|ExtrahepaticBileDuct|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C239-C241,C248-C249|ExtrahepaticBileDuct|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C239-C241,C248-C249|ExtrahepaticBileDuct|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C239-C241,C248-C249|ExtrahepaticBileDuct|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9812/3|null
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9813/3|null
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9814/3|null
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9817/3|null
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9818/3|null
C239-C241,C248-C249|ExtrahepaticBileDuct|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C239-C241,C248-C249|ExtrahepaticBileDuct|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C239-C241,C248-C249|ExtrahepaticBileDuct|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C239-C241,C248-C249|ExtrahepaticBileDuct|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C239-C241,C248-C249|ExtrahepaticBileDuct|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C239-C241,C248-C249|ExtrahepaticBileDuct|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C239-C241,C248-C249|ExtrahepaticBileDuct|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C239-C241,C248-C249|ExtrahepaticBileDuct|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C250-C254,C257-C259|Pancreas|801|Carcinoma|8010/2|InSituCancer
C250-C254,C257-C259|Pancreas|801|Carcinoma|8010/3|CarcinomaNOSDNE
C250-C254,C257-C259|Pancreas|801|Carcinoma|8011/3|MalignantEpithelioma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8012/3|LargeCellCarcinoma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8014/3|LargeCellCarcinoma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8015/3|GlassyCellCarcinoma
C250-C254,C257-C259|Pancreas|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C250-C254,C257-C259|Pancreas|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C250-C254,C257-C259|Pancreas|802|Carcinoma|8022/3|PleomorphicCarcinoma
C250-C254,C257-C259|Pancreas|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C250-C254,C257-C259|Pancreas|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C250-C254,C257-C259|Pancreas|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C250-C254,C257-C259|Pancreas|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C250-C254,C257-C259|Pancreas|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C250-C254,C257-C259|Pancreas|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C250-C254,C257-C259|Pancreas|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C250-C254,C257-C259|Pancreas|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C250-C254,C257-C259|Pancreas|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C250-C254,C257-C259|Pancreas|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C250-C254,C257-C259|Pancreas|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C250-C254,C257-C259|Pancreas|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C250-C254,C257-C259|Pancreas|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8140/3|Adenocarcinoma
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8148/2|IntraepithelialNeoplasia
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8150/3|PancreaticEndocrineCarcinoma
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8151/3|MalignantPancreaticInsulinoma
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8152/3|MalignantPancreaticGlucagonoma
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8153/3|MalignantGastrinoma
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8154/3|Adenocarcinoma
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8155/3|MalignantVipoma
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8156/3|MalignantSomatostatinoma
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8157/3|MalignantEnteroglucagonoma
C250-C254,C257-C259|Pancreas|815|EndocrineGlandNeoplasms|8158/3|ACTHProducingPituitaryGlandNeoplasm
C250-C254,C257-C259|Pancreas|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C250-C254,C257-C259|Pancreas|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C250-C254,C257-C259|Pancreas|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C250-C254,C257-C259|Pancreas|823|SolidCarcinoma|8230/2|InSituCancer
C250-C254,C257-C259|Pancreas|823|SolidCarcinoma|8230/3|SolidCarcinoma
C250-C254,C257-C259|Pancreas|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C250-C254,C257-C259|Pancreas|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C250-C254,C257-C259|Pancreas|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C250-C254,C257-C259|Pancreas|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C250-C254,C257-C259|Pancreas|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C250-C254,C257-C259|Pancreas|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C250-C254,C257-C259|Pancreas|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C250-C254,C257-C259|Pancreas|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C250-C254,C257-C259|Pancreas|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C250-C254,C257-C259|Pancreas|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C250-C254,C257-C259|Pancreas|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C250-C254,C257-C259|Pancreas|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C250-C254,C257-C259|Pancreas|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C250-C254,C257-C259|Pancreas|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C250-C254,C257-C259|Pancreas|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C250-C254,C257-C259|Pancreas|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C250-C254,C257-C259|Pancreas|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C250-C254,C257-C259|Pancreas|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C250-C254,C257-C259|Pancreas|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C250-C254,C257-C259|Pancreas|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C250-C254,C257-C259|Pancreas|845|PapillaryCystadenocarcinoma|8450/3|PapillaryCystadenocarcinoma
//C250-C254,C257-C259|Pancreas|845|PapillaryCystadenocarcinoma|8452/3|Carcinoma
C250-C254,C257-C259|Pancreas|845|PapillaryCystadenocarcinoma|8453/2|MucinousAdenocarcinoma
C250-C254,C257-C259|Pancreas|845|PapillaryCystadenocarcinoma|8453/3|MucinousAdenocarcinoma
C250-C254,C257-C259|Pancreas|847|MucinousCystadenocarcinoma|8470/2|MucinousCystadenocarcinoma
C250-C254,C257-C259|Pancreas|847|MucinousCystadenocarcinoma|8470/3|MucinousCystadenocarcinoma
C250-C254,C257-C259|Pancreas|847|MucinousCystadenocarcinoma|8471/3|PapillaryMucinousCystadenocarcinoma
C250-C254,C257-C259|Pancreas|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C250-C254,C257-C259|Pancreas|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C250-C254,C257-C259|Pancreas|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8500/2|DuctalBreastCarcinomaInSitu
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8500/3|InvasiveBreastCarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8501/2|Comedocarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8501/3|Comedocarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8503/2|IntraductalPapillaryBreastCarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8503/3|IntraductalPapillaryBreastCarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8504/2|IntracysticPapillaryBreastCarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8504/3|IntracysticPapillaryBreastCarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8507/2|MicropapillaryCarcinoma
C250-C254,C257-C259|Pancreas|850|DuctalCarcinoma|8508/3|SecretoryBreastCarcinoma
C250-C254,C257-C259|Pancreas|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C250-C254,C257-C259|Pancreas|851|MedullaryCarcinoma|8514/3|DesmoplasticNodularMedulloblastoma
C250-C254,C257-C259|Pancreas|852|IntraductalAndLobularCarcinoma|8521/3|InvasiveDuctalBreastCarcinoma
C250-C254,C257-C259|Pancreas|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C250-C254,C257-C259|Pancreas|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C250-C254,C257-C259|Pancreas|855|AcinarCellCarcinoma|8552/3|PancreaticAcinarCellCarcinoma
C250-C254,C257-C259|Pancreas|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C250-C254,C257-C259|Pancreas|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C250-C254,C257-C259|Pancreas|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C250-C254,C257-C259|Pancreas|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C250-C254,C257-C259|Pancreas|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C250-C254,C257-C259|Pancreas|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C250-C254,C257-C259|Pancreas|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C250-C254,C257-C259|Pancreas|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C250-C254,C257-C259|Pancreas|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8800/3|Sarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8801/3|SpindleCellSarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8802/3|GiantCellSarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8803/3|SmallCellSarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8804/3|SarcomaEpithelioid
C250-C254,C257-C259|Pancreas|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C250-C254,C257-C259|Pancreas|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C250-C254,C257-C259|Pancreas|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C250-C254,C257-C259|Pancreas|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C250-C254,C257-C259|Pancreas|889|MyomatousNeoplasm|8895/3|Myosarcoma
C250-C254,C257-C259|Pancreas|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C250-C254,C257-C259|Pancreas|897|Pancreatoblastoma|8971/3|Pancreatoblastoma
C250-C254,C257-C259|Pancreas|898|Carcinosarcoma|8980/3|Carcinosarcoma
C250-C254,C257-C259|Pancreas|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C250-C254,C257-C259|Pancreas|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C250-C254,C257-C259|Pancreas|959|Lymphoma|9590/3|Lymphoma
C250-C254,C257-C259|Pancreas|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C250-C254,C257-C259|Pancreas|959|Lymphoma|9596/3|CompositeLymphoma
C250-C254,C257-C259|Pancreas|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C250-C254,C257-C259|Pancreas|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C250-C254,C257-C259|Pancreas|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C250-C254,C257-C259|Pancreas|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C250-C254,C257-C259|Pancreas|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C250-C254,C257-C259|Pancreas|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C250-C254,C257-C259|Pancreas|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C250-C254,C257-C259|Pancreas|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C250-C254,C257-C259|Pancreas|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C250-C254,C257-C259|Pancreas|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C250-C254,C257-C259|Pancreas|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C250-C254,C257-C259|Pancreas|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C250-C254,C257-C259|Pancreas|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C250-C254,C257-C259|Pancreas|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C250-C254,C257-C259|Pancreas|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C250-C254,C257-C259|Pancreas|967|BCellLymphomas|9673/3|MantleCellLymphoma
C250-C254,C257-C259|Pancreas|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C250-C254,C257-C259|Pancreas|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C250-C254,C257-C259|Pancreas|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C250-C254,C257-C259|Pancreas|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C250-C254,C257-C259|Pancreas|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C250-C254,C257-C259|Pancreas|969|FollicularAdenoma|9690/3|LymphomaFollicular
C250-C254,C257-C259|Pancreas|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C250-C254,C257-C259|Pancreas|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C250-C254,C257-C259|Pancreas|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C250-C254,C257-C259|Pancreas|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C250-C254,C257-C259|Pancreas|970|TCellLymphoma|9701/3|SezarySyndrome
C250-C254,C257-C259|Pancreas|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C250-C254,C257-C259|Pancreas|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C250-C254,C257-C259|Pancreas|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C250-C254,C257-C259|Pancreas|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C250-C254,C257-C259|Pancreas|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C250-C254,C257-C259|Pancreas|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C250-C254,C257-C259|Pancreas|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C250-C254,C257-C259|Pancreas|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C250-C254,C257-C259|Pancreas|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C250-C254,C257-C259|Pancreas|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9731/3|Plasmacytoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C250-C254,C257-C259|Pancreas|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C250-C254,C257-C259|Pancreas|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C250-C254,C257-C259|Pancreas|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C250-C254,C257-C259|Pancreas|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C250-C254,C257-C259|Pancreas|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C250-C254,C257-C259|Pancreas|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C250-C254,C257-C259|Pancreas|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C250-C254,C257-C259|Pancreas|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C250-C254,C257-C259|Pancreas|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C250-C254,C257-C259|Pancreas|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C250-C254,C257-C259|Pancreas|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C250-C254,C257-C259|Pancreas|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9812/3|null
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9813/3|null
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9814/3|null
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9817/3|null
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9818/3|null
C250-C254,C257-C259|Pancreas|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C250-C254,C257-C259|Pancreas|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C250-C254,C257-C259|Pancreas|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C250-C254,C257-C259|Pancreas|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C250-C254,C257-C259|Pancreas|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C250-C254,C257-C259|Pancreas|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C250-C254,C257-C259|Pancreas|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C250-C254,C257-C259|Pancreas|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C260,C268-C269|EntireDigestiveOrgan|801|Carcinoma|8010/2|InSituCancer
C260,C268-C269|EntireDigestiveOrgan|801|Carcinoma|8010/3|CarcinomaNOSDNE
C260,C268-C269|EntireDigestiveOrgan|801|Carcinoma|8011/3|MalignantEpithelioma
C260,C268-C269|EntireDigestiveOrgan|801|Carcinoma|8012/3|LargeCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C260,C268-C269|EntireDigestiveOrgan|801|Carcinoma|8014/3|LargeCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|801|Carcinoma|8015/3|GlassyCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C260,C268-C269|EntireDigestiveOrgan|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C260,C268-C269|EntireDigestiveOrgan|802|Carcinoma|8022/3|PleomorphicCarcinoma
C260,C268-C269|EntireDigestiveOrgan|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C260,C268-C269|EntireDigestiveOrgan|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C260,C268-C269|EntireDigestiveOrgan|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C260,C268-C269|EntireDigestiveOrgan|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C260,C268-C269|EntireDigestiveOrgan|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C260,C268-C269|EntireDigestiveOrgan|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C260,C268-C269|EntireDigestiveOrgan|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C260,C268-C269|EntireDigestiveOrgan|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C260,C268-C269|EntireDigestiveOrgan|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C260,C268-C269|EntireDigestiveOrgan|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C260,C268-C269|EntireDigestiveOrgan|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C260,C268-C269|EntireDigestiveOrgan|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C260,C268-C269|EntireDigestiveOrgan|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C260,C268-C269|EntireDigestiveOrgan|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C260,C268-C269|EntireDigestiveOrgan|814|Adenocarcinoma|8140/3|Adenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C260,C268-C269|EntireDigestiveOrgan|815|EndocrineGlandNeoplasms|8152/3|MalignantPancreaticGlucagonoma
C260,C268-C269|EntireDigestiveOrgan|815|EndocrineGlandNeoplasms|8153/3|MalignantGastrinoma
C260,C268-C269|EntireDigestiveOrgan|815|EndocrineGlandNeoplasms|8156/3|MalignantSomatostatinoma
C260,C268-C269|EntireDigestiveOrgan|815|EndocrineGlandNeoplasms|8157/3|MalignantEnteroglucagonoma
C260,C268-C269|EntireDigestiveOrgan|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C260,C268-C269|EntireDigestiveOrgan|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C260,C268-C269|EntireDigestiveOrgan|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C260,C268-C269|EntireDigestiveOrgan|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C260,C268-C269|EntireDigestiveOrgan|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C260,C268-C269|EntireDigestiveOrgan|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|823|SolidCarcinoma|8230/2|InSituCancer
C260,C268-C269|EntireDigestiveOrgan|823|SolidCarcinoma|8230/3|SolidCarcinoma
C260,C268-C269|EntireDigestiveOrgan|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C260,C268-C269|EntireDigestiveOrgan|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C260,C268-C269|EntireDigestiveOrgan|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C260,C268-C269|EntireDigestiveOrgan|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C260,C268-C269|EntireDigestiveOrgan|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C260,C268-C269|EntireDigestiveOrgan|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C260,C268-C269|EntireDigestiveOrgan|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C260,C268-C269|EntireDigestiveOrgan|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C260,C268-C269|EntireDigestiveOrgan|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C260,C268-C269|EntireDigestiveOrgan|825|BronchioloalveolarAdenocarcinoma|8251/3|BronchioloalveolarAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C260,C268-C269|EntireDigestiveOrgan|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C260,C268-C269|EntireDigestiveOrgan|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C260,C268-C269|EntireDigestiveOrgan|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C260,C268-C269|EntireDigestiveOrgan|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C260,C268-C269|EntireDigestiveOrgan|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|838|CarcinomaEndometrioid|8380/3|CarcinomaEndometrioid
C260,C268-C269|EntireDigestiveOrgan|840|SweatGlandAdenocarcinoma|8401/3|ApocrineAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C260,C268-C269|EntireDigestiveOrgan|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|850|DuctalCarcinoma|8503/2|IntraductalPapillaryBreastCarcinoma
C260,C268-C269|EntireDigestiveOrgan|850|DuctalCarcinoma|8503/3|IntraductalPapillaryBreastCarcinoma
C260,C268-C269|EntireDigestiveOrgan|850|DuctalCarcinoma|8504/2|IntracysticPapillaryBreastCarcinoma
C260,C268-C269|EntireDigestiveOrgan|850|DuctalCarcinoma|8504/3|IntracysticPapillaryBreastCarcinoma
C260,C268-C269|EntireDigestiveOrgan|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C260,C268-C269|EntireDigestiveOrgan|852|IntraductalAndLobularCarcinoma|8521/3|InvasiveDuctalBreastCarcinoma
C260,C268-C269|EntireDigestiveOrgan|854|PagetDiseaseExtramammary|8542/3|PagetDiseaseExtramammary
C260,C268-C269|EntireDigestiveOrgan|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C260,C268-C269|EntireDigestiveOrgan|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C260,C268-C269|EntireDigestiveOrgan|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C260,C268-C269|EntireDigestiveOrgan|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C260,C268-C269|EntireDigestiveOrgan|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C260,C268-C269|EntireDigestiveOrgan|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C260,C268-C269|EntireDigestiveOrgan|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C260,C268-C269|EntireDigestiveOrgan|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C260,C268-C269|EntireDigestiveOrgan|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C260,C268-C269|EntireDigestiveOrgan|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C260,C268-C269|EntireDigestiveOrgan|869|MalignantExtraAdrenalParaganglioma|8693/3|MalignantExtraAdrenalParaganglioma
C260,C268-C269|EntireDigestiveOrgan|872|Melanoma|8720/2|Stage0SkinMelanoma
C260,C268-C269|EntireDigestiveOrgan|872|Melanoma|8720/3|Melanoma
C260,C268-C269|EntireDigestiveOrgan|872|Melanoma|8721/3|NodularMelanoma
C260,C268-C269|EntireDigestiveOrgan|872|Melanoma|8722/3|BalloonCellMelanoma
C260,C268-C269|EntireDigestiveOrgan|872|Melanoma|8723/3|RegressingMelanoma
C260,C268-C269|EntireDigestiveOrgan|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C260,C268-C269|EntireDigestiveOrgan|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C260,C268-C269|EntireDigestiveOrgan|874|Nevus|8745/3|DesmoplasticMelanoma
C260,C268-C269|EntireDigestiveOrgan|874|Nevus|8746/3|MucosalLentiginousMelanoma
C260,C268-C269|EntireDigestiveOrgan|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C260,C268-C269|EntireDigestiveOrgan|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C260,C268-C269|EntireDigestiveOrgan|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C260,C268-C269|EntireDigestiveOrgan|880|Sarcoma|8800/3|Sarcoma
C260,C268-C269|EntireDigestiveOrgan|880|Sarcoma|8801/3|SpindleCellSarcoma
C260,C268-C269|EntireDigestiveOrgan|880|Sarcoma|8802/3|GiantCellSarcoma
C260,C268-C269|EntireDigestiveOrgan|880|Sarcoma|8803/3|SmallCellSarcoma
C260,C268-C269|EntireDigestiveOrgan|880|Sarcoma|8804/3|SarcomaEpithelioid
C260,C268-C269|EntireDigestiveOrgan|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C260,C268-C269|EntireDigestiveOrgan|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C260,C268-C269|EntireDigestiveOrgan|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C260,C268-C269|EntireDigestiveOrgan|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C260,C268-C269|EntireDigestiveOrgan|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C260,C268-C269|EntireDigestiveOrgan|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C260,C268-C269|EntireDigestiveOrgan|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C260,C268-C269|EntireDigestiveOrgan|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C260,C268-C269|EntireDigestiveOrgan|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C260,C268-C269|EntireDigestiveOrgan|884|Myxosarcoma|8840/3|Myxosarcoma
C260,C268-C269|EntireDigestiveOrgan|885|Liposarcoma|8850/3|Liposarcoma
C260,C268-C269|EntireDigestiveOrgan|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C260,C268-C269|EntireDigestiveOrgan|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C260,C268-C269|EntireDigestiveOrgan|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C260,C268-C269|EntireDigestiveOrgan|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C260,C268-C269|EntireDigestiveOrgan|885|Liposarcoma|8855/3|Liposarcoma
C260,C268-C269|EntireDigestiveOrgan|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C260,C268-C269|EntireDigestiveOrgan|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C260,C268-C269|EntireDigestiveOrgan|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|889|MyomatousNeoplasm|8895/3|Myosarcoma
C260,C268-C269|EntireDigestiveOrgan|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C260,C268-C269|EntireDigestiveOrgan|893|StromalSarcoma|8935/3|StromalSarcoma
C260,C268-C269|EntireDigestiveOrgan|893|StromalSarcoma|8936/3|HighRiskGastrointestinalStromalTumor
C260,C268-C269|EntireDigestiveOrgan|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C260,C268-C269|EntireDigestiveOrgan|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C260,C268-C269|EntireDigestiveOrgan|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C260,C268-C269|EntireDigestiveOrgan|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C260,C268-C269|EntireDigestiveOrgan|898|Carcinosarcoma|8980/3|Carcinosarcoma
C260,C268-C269|EntireDigestiveOrgan|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C260,C268-C269|EntireDigestiveOrgan|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C260,C268-C269|EntireDigestiveOrgan|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C260,C268-C269|EntireDigestiveOrgan|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C260,C268-C269|EntireDigestiveOrgan|904|SynovialSarcoma|9040/3|SynovialSarcoma
C260,C268-C269|EntireDigestiveOrgan|904|SynovialSarcoma|9041/3|SpindleCellSynovialSarcoma
C260,C268-C269|EntireDigestiveOrgan|904|SynovialSarcoma|9042/3|EpithelialSynovialSarcoma
C260,C268-C269|EntireDigestiveOrgan|904|SynovialSarcoma|9043/3|BiphasicSynovialSarcoma
C260,C268-C269|EntireDigestiveOrgan|904|SynovialSarcoma|9044/3|ClearCellSarcomaOfSoftTissueC0206651
C260,C268-C269|EntireDigestiveOrgan|906|GermCellTumor|9060/3|Dysgerminoma
C260,C268-C269|EntireDigestiveOrgan|906|GermCellTumor|9064/3|Germinoma
C260,C268-C269|EntireDigestiveOrgan|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C260,C268-C269|EntireDigestiveOrgan|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C260,C268-C269|EntireDigestiveOrgan|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C260,C268-C269|EntireDigestiveOrgan|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C260,C268-C269|EntireDigestiveOrgan|908|Teratoma|9080/3|ImmatureTeratoma
C260,C268-C269|EntireDigestiveOrgan|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C260,C268-C269|EntireDigestiveOrgan|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C260,C268-C269|EntireDigestiveOrgan|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C260,C268-C269|EntireDigestiveOrgan|908|Teratoma|9084/3|Teratoma
C260,C268-C269|EntireDigestiveOrgan|908|Teratoma|9085/3|MixedGermCellTumor
C260,C268-C269|EntireDigestiveOrgan|910|Choriocarcinoma|9100/3|Choriocarcinoma
C260,C268-C269|EntireDigestiveOrgan|910|Choriocarcinoma|9101/3|Choriocarcinoma
C260,C268-C269|EntireDigestiveOrgan|910|Choriocarcinoma|9105/3|EpithelioidTrophoblasticTumor
C260,C268-C269|EntireDigestiveOrgan|911|Mesonephroma|9110/3|Mesonephroma
C260,C268-C269|EntireDigestiveOrgan|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C260,C268-C269|EntireDigestiveOrgan|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C260,C268-C269|EntireDigestiveOrgan|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C260,C268-C269|EntireDigestiveOrgan|914|KaposiSarcoma|9140/3|KaposiSarcoma
C260,C268-C269|EntireDigestiveOrgan|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C260,C268-C269|EntireDigestiveOrgan|917|Lymphangiosarcoma|9170/3|Lymphangiosarcoma
C260,C268-C269|EntireDigestiveOrgan|925|BoneNeoplasm|9251/3|GiantCellTumorOfSoftTissue
C260,C268-C269|EntireDigestiveOrgan|925|BoneNeoplasm|9252/3|MalignantTenosynovialGiantCellTumor
C260,C268-C269|EntireDigestiveOrgan|937|Chordoma|9370/3|Chordoma
C260,C268-C269|EntireDigestiveOrgan|937|Chordoma|9371/3|ChondroidChordoma
C260,C268-C269|EntireDigestiveOrgan|937|Chordoma|9372/3|DedifferentiatedChordoma
C260,C268-C269|EntireDigestiveOrgan|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C260,C268-C269|EntireDigestiveOrgan|950|Neuroblastoma|9500/3|Neuroblastoma
C260,C268-C269|EntireDigestiveOrgan|950|Neuroblastoma|9501/3|Medulloepithelioma
C260,C268-C269|EntireDigestiveOrgan|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C260,C268-C269|EntireDigestiveOrgan|950|Neuroblastoma|9503/3|Neuroepithelioma
C260,C268-C269|EntireDigestiveOrgan|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C260,C268-C269|EntireDigestiveOrgan|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C260,C268-C269|EntireDigestiveOrgan|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C260,C268-C269|EntireDigestiveOrgan|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C260,C268-C269|EntireDigestiveOrgan|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C260,C268-C269|EntireDigestiveOrgan|957|Perineurioma|9571/3|MalignantPerineurioma
C260,C268-C269|EntireDigestiveOrgan|959|Lymphoma|9590/3|Lymphoma
C260,C268-C269|EntireDigestiveOrgan|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C260,C268-C269|EntireDigestiveOrgan|959|Lymphoma|9596/3|CompositeLymphoma
C260,C268-C269|EntireDigestiveOrgan|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C260,C268-C269|EntireDigestiveOrgan|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C260,C268-C269|EntireDigestiveOrgan|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C260,C268-C269|EntireDigestiveOrgan|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C260,C268-C269|EntireDigestiveOrgan|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C260,C268-C269|EntireDigestiveOrgan|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C260,C268-C269|EntireDigestiveOrgan|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C260,C268-C269|EntireDigestiveOrgan|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C260,C268-C269|EntireDigestiveOrgan|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C260,C268-C269|EntireDigestiveOrgan|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C260,C268-C269|EntireDigestiveOrgan|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C260,C268-C269|EntireDigestiveOrgan|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C260,C268-C269|EntireDigestiveOrgan|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C260,C268-C269|EntireDigestiveOrgan|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C260,C268-C269|EntireDigestiveOrgan|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C260,C268-C269|EntireDigestiveOrgan|967|BCellLymphomas|9673/3|MantleCellLymphoma
C260,C268-C269|EntireDigestiveOrgan|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C260,C268-C269|EntireDigestiveOrgan|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C260,C268-C269|EntireDigestiveOrgan|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C260,C268-C269|EntireDigestiveOrgan|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C260,C268-C269|EntireDigestiveOrgan|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C260,C268-C269|EntireDigestiveOrgan|969|FollicularAdenoma|9690/3|LymphomaFollicular
C260,C268-C269|EntireDigestiveOrgan|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C260,C268-C269|EntireDigestiveOrgan|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C260,C268-C269|EntireDigestiveOrgan|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C260,C268-C269|EntireDigestiveOrgan|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C260,C268-C269|EntireDigestiveOrgan|970|TCellLymphoma|9701/3|SezarySyndrome
C260,C268-C269|EntireDigestiveOrgan|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C260,C268-C269|EntireDigestiveOrgan|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C260,C268-C269|EntireDigestiveOrgan|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C260,C268-C269|EntireDigestiveOrgan|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C260,C268-C269|EntireDigestiveOrgan|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C260,C268-C269|EntireDigestiveOrgan|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C260,C268-C269|EntireDigestiveOrgan|971|AdultNonHodgkinLymphoma|9717/3|IntestinalTCellLymphomaNOS
C260,C268-C269|EntireDigestiveOrgan|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C260,C268-C269|EntireDigestiveOrgan|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C260,C268-C269|EntireDigestiveOrgan|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C260,C268-C269|EntireDigestiveOrgan|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C260,C268-C269|EntireDigestiveOrgan|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C260,C268-C269|EntireDigestiveOrgan|973|Plasmacytoma|9731/3|Plasmacytoma
C260,C268-C269|EntireDigestiveOrgan|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C260,C268-C269|EntireDigestiveOrgan|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C260,C268-C269|EntireDigestiveOrgan|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C260,C268-C269|EntireDigestiveOrgan|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C260,C268-C269|EntireDigestiveOrgan|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C260,C268-C269|EntireDigestiveOrgan|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C260,C268-C269|EntireDigestiveOrgan|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C260,C268-C269|EntireDigestiveOrgan|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C260,C268-C269|EntireDigestiveOrgan|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C260,C268-C269|EntireDigestiveOrgan|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C260,C268-C269|EntireDigestiveOrgan|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C260,C268-C269|EntireDigestiveOrgan|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C260,C268-C269|EntireDigestiveOrgan|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C260,C268-C269|EntireDigestiveOrgan|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C260,C268-C269|EntireDigestiveOrgan|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C260,C268-C269|EntireDigestiveOrgan|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9812/3|null
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9813/3|null
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9814/3|null
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9817/3|null
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9818/3|null
C260,C268-C269|EntireDigestiveOrgan|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C260,C268-C269|EntireDigestiveOrgan|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C260,C268-C269|EntireDigestiveOrgan|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C260,C268-C269|EntireDigestiveOrgan|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C260,C268-C269|EntireDigestiveOrgan|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C260,C268-C269|EntireDigestiveOrgan|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C260,C268-C269|EntireDigestiveOrgan|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C260,C268-C269|EntireDigestiveOrgan|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C300|NasalCartilage|801|Carcinoma|8010/2|InSituCancer
C300|NasalCartilage|801|Carcinoma|8010/3|CarcinomaNOSDNE
C300|NasalCartilage|801|Carcinoma|8011/3|MalignantEpithelioma
C300|NasalCartilage|801|Carcinoma|8012/3|LargeCellCarcinoma
C300|NasalCartilage|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C300|NasalCartilage|801|Carcinoma|8014/3|LargeCellCarcinoma
C300|NasalCartilage|801|Carcinoma|8015/3|GlassyCellCarcinoma
C300|NasalCartilage|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C300|NasalCartilage|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C300|NasalCartilage|802|Carcinoma|8022/3|PleomorphicCarcinoma
C300|NasalCartilage|802|Carcinoma|8023/3|NUTCarcinoma
C300|NasalCartilage|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C300|NasalCartilage|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C300|NasalCartilage|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C300|NasalCartilage|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C300|NasalCartilage|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C300|NasalCartilage|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C300|NasalCartilage|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C300|NasalCartilage|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C300|NasalCartilage|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C300|NasalCartilage|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C300|NasalCartilage|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C300|NasalCartilage|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C300|NasalCartilage|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C300|NasalCartilage|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C300|NasalCartilage|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C300|NasalCartilage|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C300|NasalCartilage|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C300|NasalCartilage|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C300|NasalCartilage|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C300|NasalCartilage|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C300|NasalCartilage|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C300|NasalCartilage|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C300|NasalCartilage|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C300|NasalCartilage|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C300|NasalCartilage|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C300|NasalCartilage|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C300|NasalCartilage|814|Adenocarcinoma|8140/3|Adenocarcinoma
C300|NasalCartilage|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C300|NasalCartilage|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C300|NasalCartilage|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C300|NasalCartilage|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C300|NasalCartilage|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C300|NasalCartilage|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C300|NasalCartilage|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C300|NasalCartilage|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C300|NasalCartilage|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C300|NasalCartilage|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C300|NasalCartilage|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C300|NasalCartilage|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C300|NasalCartilage|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C300|NasalCartilage|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C300|NasalCartilage|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C300|NasalCartilage|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C300|NasalCartilage|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C300|NasalCartilage|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C300|NasalCartilage|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C300|NasalCartilage|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C300|NasalCartilage|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C300|NasalCartilage|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C300|NasalCartilage|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C300|NasalCartilage|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C300|NasalCartilage|872|Melanoma|8720/2|Stage0SkinMelanoma
C300|NasalCartilage|872|Melanoma|8720/3|Melanoma
C300|NasalCartilage|872|Melanoma|8721/3|NodularMelanoma
C300|NasalCartilage|872|Melanoma|8722/3|BalloonCellMelanoma
C300|NasalCartilage|872|Melanoma|8723/3|RegressingMelanoma
C300|NasalCartilage|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C300|NasalCartilage|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C300|NasalCartilage|874|Nevus|8745/3|DesmoplasticMelanoma
C300|NasalCartilage|874|Nevus|8746/3|MucosalLentiginousMelanoma
C300|NasalCartilage|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C300|NasalCartilage|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C300|NasalCartilage|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C300|NasalCartilage|880|Sarcoma|8800/3|Sarcoma
C300|NasalCartilage|880|Sarcoma|8801/3|SpindleCellSarcoma
C300|NasalCartilage|880|Sarcoma|8802/3|GiantCellSarcoma
C300|NasalCartilage|880|Sarcoma|8803/3|SmallCellSarcoma
C300|NasalCartilage|880|Sarcoma|8804/3|SarcomaEpithelioid
C300|NasalCartilage|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C300|NasalCartilage|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C300|NasalCartilage|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C300|NasalCartilage|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C300|NasalCartilage|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C300|NasalCartilage|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C300|NasalCartilage|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C300|NasalCartilage|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C300|NasalCartilage|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C300|NasalCartilage|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C300|NasalCartilage|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C300|NasalCartilage|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C300|NasalCartilage|889|MyomatousNeoplasm|8895/3|Myosarcoma
C300|NasalCartilage|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C300|NasalCartilage|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C300|NasalCartilage|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C300|NasalCartilage|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C300|NasalCartilage|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C300|NasalCartilage|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C300|NasalCartilage|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C300|NasalCartilage|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C300|NasalCartilage|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C300|NasalCartilage|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C300|NasalCartilage|904|SynovialSarcoma|9045/3|Sarcoma
C300|NasalCartilage|922|Chondrosarcoma|9220/3|Chondrosarcoma
C300|NasalCartilage|922|Chondrosarcoma|9221/3|PeriostealChondrosarcoma
C300|NasalCartilage|937|Chordoma|9370/3|Chordoma
C300|NasalCartilage|937|Chordoma|9371/3|ChondroidChordoma
C300|NasalCartilage|937|Chordoma|9372/3|DedifferentiatedChordoma
C300|NasalCartilage|950|Neuroblastoma|9500/3|Neuroblastoma
C300|NasalCartilage|950|Neuroblastoma|9501/3|Medulloepithelioma
C300|NasalCartilage|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C300|NasalCartilage|950|Neuroblastoma|9503/3|Neuroepithelioma
C300|NasalCartilage|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C300|NasalCartilage|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C300|NasalCartilage|952|OlfactoryNeurocytoma|9521/3|OlfactoryNeurocytoma
C300|NasalCartilage|952|OlfactoryNeurocytoma|9522/3|OlfactoryNeuroblastoma
C300|NasalCartilage|952|OlfactoryNeurocytoma|9523/3|OlfactoryNeuroblastoma
C300|NasalCartilage|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C300|NasalCartilage|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C300|NasalCartilage|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C300|NasalCartilage|959|Lymphoma|9590/3|Lymphoma
C300|NasalCartilage|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C300|NasalCartilage|959|Lymphoma|9596/3|CompositeLymphoma
C300|NasalCartilage|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C300|NasalCartilage|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C300|NasalCartilage|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C300|NasalCartilage|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C300|NasalCartilage|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C300|NasalCartilage|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C300|NasalCartilage|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C300|NasalCartilage|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C300|NasalCartilage|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C300|NasalCartilage|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C300|NasalCartilage|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C300|NasalCartilage|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C300|NasalCartilage|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C300|NasalCartilage|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C300|NasalCartilage|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C300|NasalCartilage|967|BCellLymphomas|9673/3|MantleCellLymphoma
C300|NasalCartilage|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C300|NasalCartilage|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C300|NasalCartilage|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C300|NasalCartilage|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C300|NasalCartilage|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C300|NasalCartilage|969|FollicularAdenoma|9690/3|LymphomaFollicular
C300|NasalCartilage|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C300|NasalCartilage|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C300|NasalCartilage|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C300|NasalCartilage|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C300|NasalCartilage|970|TCellLymphoma|9701/3|SezarySyndrome
C300|NasalCartilage|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C300|NasalCartilage|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C300|NasalCartilage|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C300|NasalCartilage|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C300|NasalCartilage|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C300|NasalCartilage|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C300|NasalCartilage|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C300|NasalCartilage|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C300|NasalCartilage|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C300|NasalCartilage|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C300|NasalCartilage|973|Plasmacytoma|9731/3|Plasmacytoma
C300|NasalCartilage|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C300|NasalCartilage|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C300|NasalCartilage|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C300|NasalCartilage|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C300|NasalCartilage|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C300|NasalCartilage|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C300|NasalCartilage|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C300|NasalCartilage|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C300|NasalCartilage|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C300|NasalCartilage|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C300|NasalCartilage|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C300|NasalCartilage|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C300|NasalCartilage|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C300|NasalCartilage|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C300|NasalCartilage|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C300|NasalCartilage|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9812/3|null
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9813/3|null
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9814/3|null
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9817/3|null
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9818/3|null
C300|NasalCartilage|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C300|NasalCartilage|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C300|NasalCartilage|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C300|NasalCartilage|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C300|NasalCartilage|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C300|NasalCartilage|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C300|NasalCartilage|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C300|NasalCartilage|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C301|MiddleEar|801|Carcinoma|8010/2|InSituCancer
C301|MiddleEar|801|Carcinoma|8010/3|CarcinomaNOSDNE
C301|MiddleEar|801|Carcinoma|8011/3|MalignantEpithelioma
C301|MiddleEar|801|Carcinoma|8012/3|LargeCellCarcinoma
C301|MiddleEar|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C301|MiddleEar|801|Carcinoma|8014/3|LargeCellCarcinoma
C301|MiddleEar|801|Carcinoma|8015/3|GlassyCellCarcinoma
C301|MiddleEar|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C301|MiddleEar|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C301|MiddleEar|802|Carcinoma|8022/3|PleomorphicCarcinoma
C301|MiddleEar|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C301|MiddleEar|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C301|MiddleEar|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C301|MiddleEar|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C301|MiddleEar|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C301|MiddleEar|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C301|MiddleEar|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C301|MiddleEar|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C301|MiddleEar|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C301|MiddleEar|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C301|MiddleEar|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C301|MiddleEar|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C301|MiddleEar|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C301|MiddleEar|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C301|MiddleEar|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C301|MiddleEar|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C301|MiddleEar|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C301|MiddleEar|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C301|MiddleEar|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C301|MiddleEar|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C301|MiddleEar|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C301|MiddleEar|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C301|MiddleEar|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C301|MiddleEar|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C301|MiddleEar|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C301|MiddleEar|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C301|MiddleEar|814|Adenocarcinoma|8140/3|Adenocarcinoma
C301|MiddleEar|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C301|MiddleEar|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C301|MiddleEar|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C301|MiddleEar|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C301|MiddleEar|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C301|MiddleEar|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C301|MiddleEar|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C301|MiddleEar|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C301|MiddleEar|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C301|MiddleEar|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C301|MiddleEar|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C301|MiddleEar|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C301|MiddleEar|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C301|MiddleEar|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C301|MiddleEar|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C301|MiddleEar|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C301|MiddleEar|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C301|MiddleEar|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C301|MiddleEar|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C301|MiddleEar|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C301|MiddleEar|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C301|MiddleEar|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C301|MiddleEar|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C301|MiddleEar|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C301|MiddleEar|872|Melanoma|8720/2|Stage0SkinMelanoma
C301|MiddleEar|872|Melanoma|8720/3|Melanoma
C301|MiddleEar|872|Melanoma|8721/3|NodularMelanoma
C301|MiddleEar|872|Melanoma|8722/3|BalloonCellMelanoma
C301|MiddleEar|872|Melanoma|8723/3|RegressingMelanoma
C301|MiddleEar|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C301|MiddleEar|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C301|MiddleEar|874|Nevus|8745/3|DesmoplasticMelanoma
C301|MiddleEar|874|Nevus|8746/3|MucosalLentiginousMelanoma
C301|MiddleEar|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C301|MiddleEar|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C301|MiddleEar|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C301|MiddleEar|880|Sarcoma|8800/3|Sarcoma
C301|MiddleEar|880|Sarcoma|8801/3|SpindleCellSarcoma
C301|MiddleEar|880|Sarcoma|8802/3|GiantCellSarcoma
C301|MiddleEar|880|Sarcoma|8803/3|SmallCellSarcoma
C301|MiddleEar|880|Sarcoma|8804/3|SarcomaEpithelioid
C301|MiddleEar|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C301|MiddleEar|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C301|MiddleEar|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C301|MiddleEar|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C301|MiddleEar|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C301|MiddleEar|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C301|MiddleEar|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C301|MiddleEar|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C301|MiddleEar|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C301|MiddleEar|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C301|MiddleEar|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C301|MiddleEar|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C301|MiddleEar|889|MyomatousNeoplasm|8895/3|Myosarcoma
C301|MiddleEar|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C301|MiddleEar|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C301|MiddleEar|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C301|MiddleEar|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C301|MiddleEar|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C301|MiddleEar|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C301|MiddleEar|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C301|MiddleEar|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C301|MiddleEar|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C301|MiddleEar|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C301|MiddleEar|937|Chordoma|9370/3|Chordoma
C301|MiddleEar|937|Chordoma|9371/3|ChondroidChordoma
C301|MiddleEar|937|Chordoma|9372/3|DedifferentiatedChordoma
C301|MiddleEar|950|Neuroblastoma|9500/3|Neuroblastoma
C301|MiddleEar|950|Neuroblastoma|9501/3|Medulloepithelioma
C301|MiddleEar|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C301|MiddleEar|950|Neuroblastoma|9503/3|Neuroepithelioma
C301|MiddleEar|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C301|MiddleEar|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C301|MiddleEar|952|OlfactoryNeurocytoma|9521/3|OlfactoryNeurocytoma
C301|MiddleEar|952|OlfactoryNeurocytoma|9522/3|OlfactoryNeuroblastoma
C301|MiddleEar|952|OlfactoryNeurocytoma|9523/3|OlfactoryNeuroblastoma
C301|MiddleEar|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C301|MiddleEar|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C301|MiddleEar|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C301|MiddleEar|957|Perineurioma|9571/3|MalignantPerineurioma
C301|MiddleEar|959|Lymphoma|9590/3|Lymphoma
C301|MiddleEar|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C301|MiddleEar|959|Lymphoma|9596/3|CompositeLymphoma
C301|MiddleEar|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C301|MiddleEar|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C301|MiddleEar|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C301|MiddleEar|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C301|MiddleEar|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C301|MiddleEar|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C301|MiddleEar|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C301|MiddleEar|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C301|MiddleEar|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C301|MiddleEar|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C301|MiddleEar|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C301|MiddleEar|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C301|MiddleEar|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C301|MiddleEar|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C301|MiddleEar|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C301|MiddleEar|967|BCellLymphomas|9673/3|MantleCellLymphoma
C301|MiddleEar|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C301|MiddleEar|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C301|MiddleEar|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C301|MiddleEar|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C301|MiddleEar|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C301|MiddleEar|969|FollicularAdenoma|9690/3|LymphomaFollicular
C301|MiddleEar|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C301|MiddleEar|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C301|MiddleEar|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C301|MiddleEar|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C301|MiddleEar|970|TCellLymphoma|9701/3|SezarySyndrome
C301|MiddleEar|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C301|MiddleEar|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C301|MiddleEar|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C301|MiddleEar|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C301|MiddleEar|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C301|MiddleEar|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C301|MiddleEar|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C301|MiddleEar|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C301|MiddleEar|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C301|MiddleEar|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C301|MiddleEar|973|Plasmacytoma|9731/3|Plasmacytoma
C301|MiddleEar|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C301|MiddleEar|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C301|MiddleEar|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C301|MiddleEar|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C301|MiddleEar|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C301|MiddleEar|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C301|MiddleEar|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C301|MiddleEar|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C301|MiddleEar|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C301|MiddleEar|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C301|MiddleEar|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C301|MiddleEar|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C301|MiddleEar|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C301|MiddleEar|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C301|MiddleEar|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C301|MiddleEar|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9812/3|null
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9813/3|null
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9814/3|null
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9817/3|null
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9818/3|null
C301|MiddleEar|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C301|MiddleEar|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C301|MiddleEar|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C301|MiddleEar|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C301|MiddleEar|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C301|MiddleEar|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C301|MiddleEar|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C301|MiddleEar|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C310-C313, C318|NasalSinus|801|Carcinoma|8010/2|InSituCancer
C310-C313, C318|NasalSinus|801|Carcinoma|8010/3|CarcinomaNOSDNE
C310-C313, C318|NasalSinus|801|Carcinoma|8011/3|MalignantEpithelioma
C310-C313, C318|NasalSinus|801|Carcinoma|8012/3|LargeCellCarcinoma
C310-C313, C318|NasalSinus|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C310-C313, C318|NasalSinus|801|Carcinoma|8014/3|LargeCellCarcinoma
C310-C313, C318|NasalSinus|801|Carcinoma|8015/3|GlassyCellCarcinoma
C310-C313, C318|NasalSinus|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C310-C313, C318|NasalSinus|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C310-C313, C318|NasalSinus|802|Carcinoma|8022/3|PleomorphicCarcinoma
C310-C313, C318|NasalSinus|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C310-C313, C318|NasalSinus|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C310-C313, C318|NasalSinus|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C310-C313, C318|NasalSinus|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C310-C313, C318|NasalSinus|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C310-C313, C318|NasalSinus|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C310-C313, C318|NasalSinus|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C310-C313, C318|NasalSinus|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C310-C313, C318|NasalSinus|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C310-C313, C318|NasalSinus|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C310-C313, C318|NasalSinus|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C310-C313, C318|NasalSinus|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C310-C313, C318|NasalSinus|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C310-C313, C318|NasalSinus|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C310-C313, C318|NasalSinus|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C310-C313, C318|NasalSinus|808|LymphoepithelialCarcinoma|8085/3|SquamousCellCarcinoma
C310-C313, C318|NasalSinus|808|LymphoepithelialCarcinoma|8086/3|SquamousCellCarcinoma
C310-C313, C318|NasalSinus|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C310-C313, C318|NasalSinus|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C310-C313, C318|NasalSinus|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C310-C313, C318|NasalSinus|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C310-C313, C318|NasalSinus|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C310-C313, C318|NasalSinus|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C310-C313, C318|NasalSinus|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C310-C313, C318|NasalSinus|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C310-C313, C318|NasalSinus|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C310-C313, C318|NasalSinus|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C310-C313, C318|NasalSinus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C310-C313, C318|NasalSinus|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C310-C313, C318|NasalSinus|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C310-C313, C318|NasalSinus|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C310-C313, C318|NasalSinus|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C310-C313, C318|NasalSinus|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C310-C313, C318|NasalSinus|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C310-C313, C318|NasalSinus|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C310-C313, C318|NasalSinus|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C310-C313, C318|NasalSinus|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C310-C313, C318|NasalSinus|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C310-C313, C318|NasalSinus|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C310-C313, C318|NasalSinus|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C310-C313, C318|NasalSinus|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C310-C313, C318|NasalSinus|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C310-C313, C318|NasalSinus|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C310-C313, C318|NasalSinus|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C310-C313, C318|NasalSinus|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C310-C313, C318|NasalSinus|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C310-C313, C318|NasalSinus|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C310-C313, C318|NasalSinus|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C310-C313, C318|NasalSinus|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C310-C313, C318|NasalSinus|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C310-C313, C318|NasalSinus|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C310-C313, C318|NasalSinus|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C310-C313, C318|NasalSinus|872|Melanoma|8720/2|Stage0SkinMelanoma
C310-C313, C318|NasalSinus|872|Melanoma|8720/3|Melanoma
C310-C313, C318|NasalSinus|872|Melanoma|8721/3|NodularMelanoma
C310-C313, C318|NasalSinus|872|Melanoma|8722/3|BalloonCellMelanoma
C310-C313, C318|NasalSinus|872|Melanoma|8723/3|RegressingMelanoma
C310-C313, C318|NasalSinus|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C310-C313, C318|NasalSinus|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C310-C313, C318|NasalSinus|874|Nevus|8745/3|DesmoplasticMelanoma
C310-C313, C318|NasalSinus|874|Nevus|8746/3|MucosalLentiginousMelanoma
C310-C313, C318|NasalSinus|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C310-C313, C318|NasalSinus|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C310-C313, C318|NasalSinus|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C310-C313, C318|NasalSinus|880|Sarcoma|8800/3|Sarcoma
C310-C313, C318|NasalSinus|880|Sarcoma|8801/3|SpindleCellSarcoma
C310-C313, C318|NasalSinus|880|Sarcoma|8802/3|GiantCellSarcoma
C310-C313, C318|NasalSinus|880|Sarcoma|8803/3|SmallCellSarcoma
C310-C313, C318|NasalSinus|880|Sarcoma|8804/3|SarcomaEpithelioid
C310-C313, C318|NasalSinus|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C310-C313, C318|NasalSinus|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C310-C313, C318|NasalSinus|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C310-C313, C318|NasalSinus|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C310-C313, C318|NasalSinus|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C310-C313, C318|NasalSinus|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C310-C313, C318|NasalSinus|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C310-C313, C318|NasalSinus|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C310-C313, C318|NasalSinus|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C310-C313, C318|NasalSinus|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C310-C313, C318|NasalSinus|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C310-C313, C318|NasalSinus|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C310-C313, C318|NasalSinus|889|MyomatousNeoplasm|8895/3|Myosarcoma
C310-C313, C318|NasalSinus|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C310-C313, C318|NasalSinus|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C310-C313, C318|NasalSinus|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C310-C313, C318|NasalSinus|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C310-C313, C318|NasalSinus|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C310-C313, C318|NasalSinus|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C310-C313, C318|NasalSinus|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C310-C313, C318|NasalSinus|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C310-C313, C318|NasalSinus|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C310-C313, C318|NasalSinus|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C310-C313, C318|NasalSinus|904|SynovialSarcoma|9045/3|Sarcoma
C310-C313, C318|NasalSinus|937|Chordoma|9370/3|Chordoma
C310-C313, C318|NasalSinus|937|Chordoma|9371/3|ChondroidChordoma
C310-C313, C318|NasalSinus|937|Chordoma|9372/3|DedifferentiatedChordoma
C310-C313, C318|NasalSinus|950|Neuroblastoma|9500/3|Neuroblastoma
C310-C313, C318|NasalSinus|950|Neuroblastoma|9501/3|Medulloepithelioma
C310-C313, C318|NasalSinus|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C310-C313, C318|NasalSinus|950|Neuroblastoma|9503/3|Neuroepithelioma
C310-C313, C318|NasalSinus|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C310-C313, C318|NasalSinus|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C310-C313, C318|NasalSinus|952|OlfactoryNeurocytoma|9521/3|OlfactoryNeurocytoma
C310-C313, C318|NasalSinus|952|OlfactoryNeurocytoma|9522/3|OlfactoryNeuroblastoma
C310-C313, C318|NasalSinus|952|OlfactoryNeurocytoma|9523/3|OlfactoryNeuroblastoma
C310-C313, C318|NasalSinus|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C310-C313, C318|NasalSinus|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C310-C313, C318|NasalSinus|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C310-C313, C318|NasalSinus|957|Perineurioma|9571/3|MalignantPerineurioma
C310-C313, C318|NasalSinus|959|Lymphoma|9590/3|Lymphoma
C310-C313, C318|NasalSinus|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C310-C313, C318|NasalSinus|959|Lymphoma|9596/3|CompositeLymphoma
C310-C313, C318|NasalSinus|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C310-C313, C318|NasalSinus|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C310-C313, C318|NasalSinus|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C310-C313, C318|NasalSinus|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C310-C313, C318|NasalSinus|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C310-C313, C318|NasalSinus|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C310-C313, C318|NasalSinus|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C310-C313, C318|NasalSinus|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C310-C313, C318|NasalSinus|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C310-C313, C318|NasalSinus|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C310-C313, C318|NasalSinus|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C310-C313, C318|NasalSinus|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C310-C313, C318|NasalSinus|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C310-C313, C318|NasalSinus|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C310-C313, C318|NasalSinus|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C310-C313, C318|NasalSinus|967|BCellLymphomas|9673/3|MantleCellLymphoma
C310-C313, C318|NasalSinus|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C310-C313, C318|NasalSinus|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C310-C313, C318|NasalSinus|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C310-C313, C318|NasalSinus|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C310-C313, C318|NasalSinus|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C310-C313, C318|NasalSinus|969|FollicularAdenoma|9690/3|LymphomaFollicular
C310-C313, C318|NasalSinus|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C310-C313, C318|NasalSinus|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C310-C313, C318|NasalSinus|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C310-C313, C318|NasalSinus|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C310-C313, C318|NasalSinus|970|TCellLymphoma|9701/3|SezarySyndrome
C310-C313, C318|NasalSinus|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C310-C313, C318|NasalSinus|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C310-C313, C318|NasalSinus|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C310-C313, C318|NasalSinus|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C310-C313, C318|NasalSinus|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C310-C313, C318|NasalSinus|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C310-C313, C318|NasalSinus|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C310-C313, C318|NasalSinus|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C310-C313, C318|NasalSinus|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C310-C313, C318|NasalSinus|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C310-C313, C318|NasalSinus|973|Plasmacytoma|9731/3|Plasmacytoma
C310-C313, C318|NasalSinus|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C310-C313, C318|NasalSinus|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C310-C313, C318|NasalSinus|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C310-C313, C318|NasalSinus|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C310-C313, C318|NasalSinus|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C310-C313, C318|NasalSinus|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C310-C313, C318|NasalSinus|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C310-C313, C318|NasalSinus|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C310-C313, C318|NasalSinus|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C310-C313, C318|NasalSinus|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C310-C313, C318|NasalSinus|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C310-C313, C318|NasalSinus|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C310-C313, C318|NasalSinus|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C310-C313, C318|NasalSinus|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C310-C313, C318|NasalSinus|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C310-C313, C318|NasalSinus|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9812/3|null
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9813/3|null
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9814/3|null
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9817/3|null
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9818/3|null
C310-C313, C318|NasalSinus|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C310-C313, C318|NasalSinus|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C310-C313, C318|NasalSinus|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C310-C313, C318|NasalSinus|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C310-C313, C318|NasalSinus|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C310-C313, C318|NasalSinus|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C310-C313, C318|NasalSinus|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C310-C313, C318|NasalSinus|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C319|NasalSinus|801|Carcinoma|8010/2|InSituCancer
C319|NasalSinus|801|Carcinoma|8010/3|CarcinomaNOSDNE
C319|NasalSinus|801|Carcinoma|8011/3|MalignantEpithelioma
C319|NasalSinus|801|Carcinoma|8012/3|LargeCellCarcinoma
C319|NasalSinus|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C319|NasalSinus|801|Carcinoma|8014/3|LargeCellCarcinoma
C319|NasalSinus|801|Carcinoma|8015/3|GlassyCellCarcinoma
C319|NasalSinus|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C319|NasalSinus|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C319|NasalSinus|802|Carcinoma|8022/3|PleomorphicCarcinoma
C319|NasalSinus|802|Carcinoma|8023/3|NUTCarcinoma
C319|NasalSinus|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C319|NasalSinus|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C319|NasalSinus|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C319|NasalSinus|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C319|NasalSinus|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C319|NasalSinus|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C319|NasalSinus|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C319|NasalSinus|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C319|NasalSinus|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C319|NasalSinus|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C319|NasalSinus|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C319|NasalSinus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C319|NasalSinus|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C319|NasalSinus|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C319|NasalSinus|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C319|NasalSinus|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C319|NasalSinus|808|LymphoepithelialCarcinoma|8085/3|SquamousCellCarcinoma
C319|NasalSinus|808|LymphoepithelialCarcinoma|8086/3|SquamousCellCarcinoma
C319|NasalSinus|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C319|NasalSinus|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C319|NasalSinus|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C319|NasalSinus|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C319|NasalSinus|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C319|NasalSinus|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C319|NasalSinus|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C319|NasalSinus|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C319|NasalSinus|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C319|NasalSinus|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C319|NasalSinus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C319|NasalSinus|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C319|NasalSinus|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C319|NasalSinus|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C319|NasalSinus|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C319|NasalSinus|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C319|NasalSinus|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C319|NasalSinus|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C319|NasalSinus|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C319|NasalSinus|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C319|NasalSinus|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C319|NasalSinus|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C319|NasalSinus|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C319|NasalSinus|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C319|NasalSinus|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C319|NasalSinus|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C319|NasalSinus|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C319|NasalSinus|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C319|NasalSinus|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C319|NasalSinus|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C319|NasalSinus|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C319|NasalSinus|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C319|NasalSinus|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C319|NasalSinus|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C319|NasalSinus|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C319|NasalSinus|872|Melanoma|8720/2|Stage0SkinMelanoma
C319|NasalSinus|872|Melanoma|8720/3|Melanoma
C319|NasalSinus|872|Melanoma|8721/3|NodularMelanoma
C319|NasalSinus|872|Melanoma|8722/3|BalloonCellMelanoma
C319|NasalSinus|872|Melanoma|8723/3|RegressingMelanoma
C319|NasalSinus|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C319|NasalSinus|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C319|NasalSinus|874|Nevus|8745/3|DesmoplasticMelanoma
C319|NasalSinus|874|Nevus|8746/3|MucosalLentiginousMelanoma
C319|NasalSinus|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C319|NasalSinus|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C319|NasalSinus|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C319|NasalSinus|880|Sarcoma|8800/3|Sarcoma
C319|NasalSinus|880|Sarcoma|8801/3|SpindleCellSarcoma
C319|NasalSinus|880|Sarcoma|8802/3|GiantCellSarcoma
C319|NasalSinus|880|Sarcoma|8803/3|SmallCellSarcoma
C319|NasalSinus|880|Sarcoma|8804/3|SarcomaEpithelioid
C319|NasalSinus|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C319|NasalSinus|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C319|NasalSinus|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C319|NasalSinus|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C319|NasalSinus|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C319|NasalSinus|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C319|NasalSinus|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C319|NasalSinus|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C319|NasalSinus|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C319|NasalSinus|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C319|NasalSinus|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C319|NasalSinus|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C319|NasalSinus|889|MyomatousNeoplasm|8895/3|Myosarcoma
C319|NasalSinus|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C319|NasalSinus|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C319|NasalSinus|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C319|NasalSinus|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C319|NasalSinus|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C319|NasalSinus|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C319|NasalSinus|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C319|NasalSinus|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C319|NasalSinus|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C319|NasalSinus|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C319|NasalSinus|904|SynovialSarcoma|9045/3|Sarcoma
C319|NasalSinus|937|Chordoma|9370/3|Chordoma
C319|NasalSinus|937|Chordoma|9371/3|ChondroidChordoma
C319|NasalSinus|937|Chordoma|9372/3|DedifferentiatedChordoma
C319|NasalSinus|950|Neuroblastoma|9500/3|Neuroblastoma
C319|NasalSinus|950|Neuroblastoma|9501/3|Medulloepithelioma
C319|NasalSinus|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C319|NasalSinus|950|Neuroblastoma|9503/3|Neuroepithelioma
C319|NasalSinus|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C319|NasalSinus|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C319|NasalSinus|952|OlfactoryNeurocytoma|9521/3|OlfactoryNeurocytoma
C319|NasalSinus|952|OlfactoryNeurocytoma|9522/3|OlfactoryNeuroblastoma
C319|NasalSinus|952|OlfactoryNeurocytoma|9523/3|OlfactoryNeuroblastoma
C319|NasalSinus|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C319|NasalSinus|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C319|NasalSinus|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C319|NasalSinus|957|Perineurioma|9571/3|MalignantPerineurioma
C319|NasalSinus|959|Lymphoma|9590/3|Lymphoma
C319|NasalSinus|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C319|NasalSinus|959|Lymphoma|9596/3|CompositeLymphoma
C319|NasalSinus|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C319|NasalSinus|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C319|NasalSinus|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C319|NasalSinus|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C319|NasalSinus|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C319|NasalSinus|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C319|NasalSinus|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C319|NasalSinus|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C319|NasalSinus|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C319|NasalSinus|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C319|NasalSinus|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C319|NasalSinus|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C319|NasalSinus|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C319|NasalSinus|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C319|NasalSinus|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C319|NasalSinus|967|BCellLymphomas|9673/3|MantleCellLymphoma
C319|NasalSinus|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C319|NasalSinus|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C319|NasalSinus|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C319|NasalSinus|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C319|NasalSinus|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C319|NasalSinus|969|FollicularAdenoma|9690/3|LymphomaFollicular
C319|NasalSinus|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C319|NasalSinus|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C319|NasalSinus|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C319|NasalSinus|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C319|NasalSinus|970|TCellLymphoma|9701/3|SezarySyndrome
C319|NasalSinus|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C319|NasalSinus|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C319|NasalSinus|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C319|NasalSinus|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C319|NasalSinus|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C319|NasalSinus|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C319|NasalSinus|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C319|NasalSinus|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C319|NasalSinus|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C319|NasalSinus|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C319|NasalSinus|973|Plasmacytoma|9731/3|Plasmacytoma
C319|NasalSinus|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C319|NasalSinus|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C319|NasalSinus|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C319|NasalSinus|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C319|NasalSinus|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C319|NasalSinus|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C319|NasalSinus|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C319|NasalSinus|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C319|NasalSinus|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C319|NasalSinus|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C319|NasalSinus|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C319|NasalSinus|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C319|NasalSinus|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C319|NasalSinus|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C319|NasalSinus|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C319|NasalSinus|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9812/3|null
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9813/3|null
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9814/3|null
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9817/3|null
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9818/3|null
C319|NasalSinus|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C319|NasalSinus|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C319|NasalSinus|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C319|NasalSinus|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C319|NasalSinus|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C319|NasalSinus|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C319|NasalSinus|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C319|NasalSinus|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C320-C323,C328-C329|Larynx|801|Carcinoma|8010/2|InSituCancer
C320-C323,C328-C329|Larynx|801|Carcinoma|8010/3|CarcinomaNOSDNE
C320-C323,C328-C329|Larynx|801|Carcinoma|8011/3|MalignantEpithelioma
C320-C323,C328-C329|Larynx|801|Carcinoma|8012/3|LargeCellCarcinoma
C320-C323,C328-C329|Larynx|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C320-C323,C328-C329|Larynx|801|Carcinoma|8014/3|LargeCellCarcinoma
C320-C323,C328-C329|Larynx|801|Carcinoma|8015/3|GlassyCellCarcinoma
C320-C323,C328-C329|Larynx|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C320-C323,C328-C329|Larynx|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C320-C323,C328-C329|Larynx|802|Carcinoma|8022/3|PleomorphicCarcinoma
C320-C323,C328-C329|Larynx|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C320-C323,C328-C329|Larynx|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C320-C323,C328-C329|Larynx|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C320-C323,C328-C329|Larynx|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C320-C323,C328-C329|Larynx|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C320-C323,C328-C329|Larynx|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C320-C323,C328-C329|Larynx|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C320-C323,C328-C329|Larynx|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C320-C323,C328-C329|Larynx|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C320-C323,C328-C329|Larynx|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C320-C323,C328-C329|Larynx|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C320-C323,C328-C329|Larynx|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C320-C323,C328-C329|Larynx|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C320-C323,C328-C329|Larynx|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C320-C323,C328-C329|Larynx|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C320-C323,C328-C329|Larynx|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C320-C323,C328-C329|Larynx|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C320-C323,C328-C329|Larynx|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C320-C323,C328-C329|Larynx|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C320-C323,C328-C329|Larynx|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C320-C323,C328-C329|Larynx|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C320-C323,C328-C329|Larynx|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C320-C323,C328-C329|Larynx|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C320-C323,C328-C329|Larynx|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C320-C323,C328-C329|Larynx|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C320-C323,C328-C329|Larynx|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C320-C323,C328-C329|Larynx|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C320-C323,C328-C329|Larynx|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C320-C323,C328-C329|Larynx|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C320-C323,C328-C329|Larynx|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C320-C323,C328-C329|Larynx|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C320-C323,C328-C329|Larynx|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C320-C323,C328-C329|Larynx|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C320-C323,C328-C329|Larynx|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C320-C323,C328-C329|Larynx|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C320-C323,C328-C329|Larynx|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C320-C323,C328-C329|Larynx|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C320-C323,C328-C329|Larynx|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C320-C323,C328-C329|Larynx|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8800/3|Sarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8801/3|SpindleCellSarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8802/3|GiantCellSarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8803/3|SmallCellSarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8804/3|SarcomaEpithelioid
C320-C323,C328-C329|Larynx|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C320-C323,C328-C329|Larynx|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C320-C323,C328-C329|Larynx|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C320-C323,C328-C329|Larynx|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C320-C323,C328-C329|Larynx|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C320-C323,C328-C329|Larynx|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C320-C323,C328-C329|Larynx|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C320-C323,C328-C329|Larynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C320-C323,C328-C329|Larynx|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C320-C323,C328-C329|Larynx|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C320-C323,C328-C329|Larynx|922|Chondrosarcoma|9220/3|Chondrosarcoma
C320-C323,C328-C329|Larynx|922|Chondrosarcoma|9221/3|PeriostealChondrosarcoma
C320-C323,C328-C329|Larynx|959|Lymphoma|9590/3|Lymphoma
C320-C323,C328-C329|Larynx|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C320-C323,C328-C329|Larynx|959|Lymphoma|9596/3|CompositeLymphoma
C320-C323,C328-C329|Larynx|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C320-C323,C328-C329|Larynx|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C320-C323,C328-C329|Larynx|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C320-C323,C328-C329|Larynx|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C320-C323,C328-C329|Larynx|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C320-C323,C328-C329|Larynx|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C320-C323,C328-C329|Larynx|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C320-C323,C328-C329|Larynx|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C320-C323,C328-C329|Larynx|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C320-C323,C328-C329|Larynx|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C320-C323,C328-C329|Larynx|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C320-C323,C328-C329|Larynx|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C320-C323,C328-C329|Larynx|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C320-C323,C328-C329|Larynx|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C320-C323,C328-C329|Larynx|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C320-C323,C328-C329|Larynx|967|BCellLymphomas|9673/3|MantleCellLymphoma
C320-C323,C328-C329|Larynx|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C320-C323,C328-C329|Larynx|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C320-C323,C328-C329|Larynx|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C320-C323,C328-C329|Larynx|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C320-C323,C328-C329|Larynx|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C320-C323,C328-C329|Larynx|969|FollicularAdenoma|9690/3|LymphomaFollicular
C320-C323,C328-C329|Larynx|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C320-C323,C328-C329|Larynx|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C320-C323,C328-C329|Larynx|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C320-C323,C328-C329|Larynx|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C320-C323,C328-C329|Larynx|970|TCellLymphoma|9701/3|SezarySyndrome
C320-C323,C328-C329|Larynx|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C320-C323,C328-C329|Larynx|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C320-C323,C328-C329|Larynx|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C320-C323,C328-C329|Larynx|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C320-C323,C328-C329|Larynx|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C320-C323,C328-C329|Larynx|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C320-C323,C328-C329|Larynx|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C320-C323,C328-C329|Larynx|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C320-C323,C328-C329|Larynx|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C320-C323,C328-C329|Larynx|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9731/3|Plasmacytoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C320-C323,C328-C329|Larynx|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C320-C323,C328-C329|Larynx|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C320-C323,C328-C329|Larynx|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C320-C323,C328-C329|Larynx|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C320-C323,C328-C329|Larynx|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C320-C323,C328-C329|Larynx|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C320-C323,C328-C329|Larynx|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C320-C323,C328-C329|Larynx|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C320-C323,C328-C329|Larynx|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C320-C323,C328-C329|Larynx|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C320-C323,C328-C329|Larynx|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C320-C323,C328-C329|Larynx|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9812/3|null
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9813/3|null
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9814/3|null
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9817/3|null
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9818/3|null
C320-C323,C328-C329|Larynx|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C320-C323,C328-C329|Larynx|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C320-C323,C328-C329|Larynx|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C320-C323,C328-C329|Larynx|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C320-C323,C328-C329|Larynx|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C320-C323,C328-C329|Larynx|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C320-C323,C328-C329|Larynx|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C320-C323,C328-C329|Larynx|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C339|Trachea|801|Carcinoma|8010/2|InSituCancer
C339|Trachea|801|Carcinoma|8010/3|CarcinomaNOSDNE
C339|Trachea|801|Carcinoma|8011/3|MalignantEpithelioma
C339|Trachea|801|Carcinoma|8012/3|LargeCellCarcinoma
C339|Trachea|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C339|Trachea|801|Carcinoma|8014/3|LargeCellCarcinoma
C339|Trachea|801|Carcinoma|8015/3|GlassyCellCarcinoma
C339|Trachea|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C339|Trachea|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C339|Trachea|802|Carcinoma|8022/3|PleomorphicCarcinoma
C339|Trachea|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C339|Trachea|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C339|Trachea|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C339|Trachea|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C339|Trachea|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C339|Trachea|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C339|Trachea|804|NonSmallCellCarcinoma|8046/3|NonSmallCellCarcinoma
C339|Trachea|804|NonSmallCellCarcinoma|8046/6|MetastaticLungCarcinoma
C339|Trachea|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C339|Trachea|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C339|Trachea|804|SmallCellCarcinoma|8042/3|OatCell
C339|Trachea|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C339|Trachea|804|SmallCellCarcinoma|8044/3|SmallCellIntermediateCellCarcinoma
C339|Trachea|804|SmallCellCarcinoma|8045/3|CombinedSmallCellLungCarcinoma
C339|Trachea|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C339|Trachea|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C339|Trachea|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C339|Trachea|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C339|Trachea|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C339|Trachea|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C339|Trachea|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C339|Trachea|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C339|Trachea|814|Adenocarcinoma|8140/3|Adenocarcinoma
C339|Trachea|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C339|Trachea|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C339|Trachea|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C339|Trachea|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C339|Trachea|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C339|Trachea|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C339|Trachea|825|BronchioloalveolarAdenocarcinoma|8250/3|LepidicPredominantAdenocarcinoma
C339|Trachea|825|BronchioloalveolarAdenocarcinoma|8252/3|NonMucinousLungAdenocarcinomaInSitu
C339|Trachea|825|BronchioloalveolarAdenocarcinoma|8253/3|MucinousAdenocarcinoma
C339|Trachea|825|BronchioloalveolarAdenocarcinoma|8254/3|MixedSubtypeAdenocarcinomaOfLung
C339|Trachea|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C339|Trachea|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C339|Trachea|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C339|Trachea|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C339|Trachea|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C339|Trachea|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C339|Trachea|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C339|Trachea|880|Sarcoma|8800/3|Sarcoma
C339|Trachea|880|Sarcoma|8801/3|SpindleCellSarcoma
C339|Trachea|880|Sarcoma|8802/3|GiantCellSarcoma
C339|Trachea|880|Sarcoma|8803/3|SmallCellSarcoma
C339|Trachea|880|Sarcoma|8804/3|SarcomaEpithelioid
C339|Trachea|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C339|Trachea|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C339|Trachea|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C339|Trachea|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C339|Trachea|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C339|Trachea|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C339|Trachea|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C339|Trachea|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C339|Trachea|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C339|Trachea|897|Hepatoblastoma|8972/3|PulmonaryBlastoma
C339|Trachea|897|Hepatoblastoma|8973/3|PleuropulmonaryBlastoma
C339|Trachea|922|Chondrosarcoma|9220/3|Chondrosarcoma
C339|Trachea|922|Chondrosarcoma|9221/3|PeriostealChondrosarcoma
C339|Trachea|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C339|Trachea|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C340-C343,C348-C349|Bronchus|801|Carcinoma|8010/2|InSituCancer
C340-C343,C348-C349|Bronchus|801|Carcinoma|8010/3|CarcinomaNOSDNE
C340-C343,C348-C349|Bronchus|801|Carcinoma|8011/3|MalignantEpithelioma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8012/3|LargeCellCarcinoma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8014/3|LargeCellCarcinoma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8015/3|GlassyCellCarcinoma
C340-C343,C348-C349|Bronchus|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C340-C343,C348-C349|Bronchus|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C340-C343,C348-C349|Bronchus|802|Carcinoma|8022/3|PleomorphicCarcinoma
C340-C343,C348-C349|Bronchus|802|Carcinoma|8023/3|NUTCarcinoma
C340-C343,C348-C349|Bronchus|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C340-C343,C348-C349|Bronchus|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C340-C343,C348-C349|Bronchus|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C340-C343,C348-C349|Bronchus|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C340-C343,C348-C349|Bronchus|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C340-C343,C348-C349|Bronchus|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C340-C343,C348-C349|Bronchus|804|NonSmallCellCarcinoma|8046/3|NonSmallCellCarcinoma
C340-C343,C348-C349|Bronchus|804|NonSmallCellCarcinoma|8046/6|MetastaticLungCarcinoma
C340-C343,C348-C349|Bronchus|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C340-C343,C348-C349|Bronchus|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C340-C343,C348-C349|Bronchus|804|SmallCellCarcinoma|8042/3|SmallCellCarcinoma
C340-C343,C348-C349|Bronchus|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C340-C343,C348-C349|Bronchus|804|SmallCellCarcinoma|8044/3|SmallCellIntermediateCellCarcinoma
C340-C343,C348-C349|Bronchus|804|SmallCellCarcinoma|8045/3|CombinedSmallCellLungCarcinoma
C340-C343,C348-C349|Bronchus|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C340-C343,C348-C349|Bronchus|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C340-C343,C348-C349|Bronchus|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C340-C343,C348-C349|Bronchus|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C340-C343,C348-C349|Bronchus|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C340-C343,C348-C349|Bronchus|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C340-C343,C348-C349|Bronchus|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C340-C343,C348-C349|Bronchus|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C340-C343,C348-C349|Bronchus|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C340-C343,C348-C349|Bronchus|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8140/1|LungCarcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C340-C343,C348-C349|Bronchus|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C340-C343,C348-C349|Bronchus|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C340-C343,C348-C349|Bronchus|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C340-C343,C348-C349|Bronchus|823|SolidCarcinoma|8230/2|InSituCancer
C340-C343,C348-C349|Bronchus|823|SolidCarcinoma|8230/3|SolidCarcinoma
C340-C343,C348-C349|Bronchus|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C340-C343,C348-C349|Bronchus|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C340-C343,C348-C349|Bronchus|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C340-C343,C348-C349|Bronchus|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C340-C343,C348-C349|Bronchus|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C340-C343,C348-C349|Bronchus|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C340-C343,C348-C349|Bronchus|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C340-C343,C348-C349|Bronchus|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C340-C343,C348-C349|Bronchus|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8250/2|NonmucinousAdenocarcinomaInSitu
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8250/3|LepidicPredominantAdenocarcinoma
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8251/3|BronchioloalveolarAdenocarcinoma
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8252/3|NonMucinousLungAdenocarcinomaInSitu
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8253/2|MucinousAdenocarcinomaInSitu
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8253/3|MucinousAdenocarcinoma
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8254/3|MixedSubtypeAdenocarcinomaOfLung
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8256/3|InvasiveMucinousLungAdenocarcinoma
C340-C343,C348-C349|Bronchus|825|BronchioloalveolarAdenocarcinoma|8257/3|MucinousAdenocarcinoma
C340-C343,C348-C349|Bronchus|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C340-C343,C348-C349|Bronchus|826|PapillaryAdenocarcinoma|8265/3|MicropapillaryCarcinoma
C340-C343,C348-C349|Bronchus|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C340-C343,C348-C349|Bronchus|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C340-C343,C348-C349|Bronchus|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C340-C343,C348-C349|Bronchus|833|FollicularThyroidCarcinoma|8333/3|FetalAdenocarcinoma
C340-C343,C348-C349|Bronchus|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C340-C343,C348-C349|Bronchus|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C340-C343,C348-C349|Bronchus|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C340-C343,C348-C349|Bronchus|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C340-C343,C348-C349|Bronchus|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C340-C343,C348-C349|Bronchus|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C340-C343,C348-C349|Bronchus|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C340-C343,C348-C349|Bronchus|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C340-C343,C348-C349|Bronchus|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C340-C343,C348-C349|Bronchus|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C340-C343,C348-C349|Bronchus|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C340-C343,C348-C349|Bronchus|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C340-C343,C348-C349|Bronchus|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C340-C343,C348-C349|Bronchus|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C340-C343,C348-C349|Bronchus|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C340-C343,C348-C349|Bronchus|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C340-C343,C348-C349|Bronchus|871|MalignantGlomusTumor|8714/3|MalignantPEComa
C340-C343,C348-C349|Bronchus|880|Sarcoma|8800/3|Sarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8801/3|SpindleCellSarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8802/3|GiantCellSarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8803/3|SmallCellSarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8804/3|SarcomaEpithelioid
C340-C343,C348-C349|Bronchus|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C340-C343,C348-C349|Bronchus|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C340-C343,C348-C349|Bronchus|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C340-C343,C348-C349|Bronchus|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C340-C343,C348-C349|Bronchus|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C340-C343,C348-C349|Bronchus|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C340-C343,C348-C349|Bronchus|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C340-C343,C348-C349|Bronchus|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C340-C343,C348-C349|Bronchus|884|Myxosarcoma|8842/3|Sarcoma
C340-C343,C348-C349|Bronchus|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C340-C343,C348-C349|Bronchus|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C340-C343,C348-C349|Bronchus|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C340-C343,C348-C349|Bronchus|889|MyomatousNeoplasm|8895/3|Myosarcoma
C340-C343,C348-C349|Bronchus|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C340-C343,C348-C349|Bronchus|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C340-C343,C348-C349|Bronchus|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C340-C343,C348-C349|Bronchus|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C340-C343,C348-C349|Bronchus|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C340-C343,C348-C349|Bronchus|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C340-C343,C348-C349|Bronchus|897|Hepatoblastoma|8972/3|PulmonaryBlastoma
C340-C343,C348-C349|Bronchus|897|Hepatoblastoma|8973/3|PleuropulmonaryBlastoma
C340-C343,C348-C349|Bronchus|898|Carcinosarcoma|8980/3|Carcinosarcoma
C340-C343,C348-C349|Bronchus|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C340-C343,C348-C349|Bronchus|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C340-C343,C348-C349|Bronchus|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C340-C343,C348-C349|Bronchus|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C340-C343,C348-C349|Bronchus|905|MalignantMesothelioma|9050/3|MalignantMesothelioma
C340-C343,C348-C349|Bronchus|905|MalignantMesothelioma|9051/3|SarcomatoidMesothelioma
C340-C343,C348-C349|Bronchus|905|MalignantMesothelioma|9052/3|Mesothelioma
C340-C343,C348-C349|Bronchus|905|MalignantMesothelioma|9053/3|BiphasicMesothelioma
C340-C343,C348-C349|Bronchus|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C340-C343,C348-C349|Bronchus|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C340-C343,C348-C349|Bronchus|913|Hemangioendothelioma|9137/3|IntimalSarcoma
C340-C343,C348-C349|Bronchus|914|KaposiSarcoma|9140/3|KaposiSarcoma
C340-C343,C348-C349|Bronchus|959|Lymphoma|9590/3|Lymphoma
C340-C343,C348-C349|Bronchus|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C340-C343,C348-C349|Bronchus|959|Lymphoma|9596/3|CompositeLymphoma
C340-C343,C348-C349|Bronchus|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C340-C343,C348-C349|Bronchus|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C340-C343,C348-C349|Bronchus|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C340-C343,C348-C349|Bronchus|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C340-C343,C348-C349|Bronchus|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C340-C343,C348-C349|Bronchus|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C340-C343,C348-C349|Bronchus|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C340-C343,C348-C349|Bronchus|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C340-C343,C348-C349|Bronchus|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C340-C343,C348-C349|Bronchus|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C340-C343,C348-C349|Bronchus|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C340-C343,C348-C349|Bronchus|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C340-C343,C348-C349|Bronchus|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C340-C343,C348-C349|Bronchus|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C340-C343,C348-C349|Bronchus|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C340-C343,C348-C349|Bronchus|967|BCellLymphomas|9673/3|MantleCellLymphoma
C340-C343,C348-C349|Bronchus|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C340-C343,C348-C349|Bronchus|967|BCellLymphomas|9678/3|PrimaryEffusionLymphoma
C340-C343,C348-C349|Bronchus|967|BCellLymphomas|9679/3|MediastinalLargeBcellLymphoma
C340-C343,C348-C349|Bronchus|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C340-C343,C348-C349|Bronchus|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C340-C343,C348-C349|Bronchus|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C340-C343,C348-C349|Bronchus|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C340-C343,C348-C349|Bronchus|969|FollicularAdenoma|9690/3|LymphomaFollicular
C340-C343,C348-C349|Bronchus|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C340-C343,C348-C349|Bronchus|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C340-C343,C348-C349|Bronchus|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C340-C343,C348-C349|Bronchus|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C340-C343,C348-C349|Bronchus|970|TCellLymphoma|9701/3|SezarySyndrome
C340-C343,C348-C349|Bronchus|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C340-C343,C348-C349|Bronchus|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C340-C343,C348-C349|Bronchus|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C340-C343,C348-C349|Bronchus|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C340-C343,C348-C349|Bronchus|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C340-C343,C348-C349|Bronchus|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C340-C343,C348-C349|Bronchus|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C340-C343,C348-C349|Bronchus|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C340-C343,C348-C349|Bronchus|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C340-C343,C348-C349|Bronchus|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9731/3|Plasmacytoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C340-C343,C348-C349|Bronchus|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C340-C343,C348-C349|Bronchus|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C340-C343,C348-C349|Bronchus|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C340-C343,C348-C349|Bronchus|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C340-C343,C348-C349|Bronchus|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C340-C343,C348-C349|Bronchus|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C340-C343,C348-C349|Bronchus|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C340-C343,C348-C349|Bronchus|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C340-C343,C348-C349|Bronchus|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C340-C343,C348-C349|Bronchus|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C340-C343,C348-C349|Bronchus|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C340-C343,C348-C349|Bronchus|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9812/3|null
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9813/3|null
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9814/3|null
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9817/3|null
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9818/3|null
C340-C343,C348-C349|Bronchus|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C340-C343,C348-C349|Bronchus|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C340-C343,C348-C349|Bronchus|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C340-C343,C348-C349|Bronchus|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C340-C343,C348-C349|Bronchus|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C340-C343,C348-C349|Bronchus|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C340-C343,C348-C349|Bronchus|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C340-C343,C348-C349|Bronchus|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C379|ThymusGland|801|Carcinoma|8010/2|InSituCancer
C379|ThymusGland|801|Carcinoma|8010/3|CarcinomaNOSDNE
C379|ThymusGland|801|Carcinoma|8011/3|MalignantEpithelioma
C379|ThymusGland|801|Carcinoma|8012/3|LargeCellCarcinoma
C379|ThymusGland|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C379|ThymusGland|801|Carcinoma|8014/3|LargeCellCarcinoma
C379|ThymusGland|801|Carcinoma|8015/3|GlassyCellCarcinoma
C379|ThymusGland|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C379|ThymusGland|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C379|ThymusGland|802|Carcinoma|8022/3|PleomorphicCarcinoma
C379|ThymusGland|802|Carcinoma|8023/3|NUTCarcinoma
C379|ThymusGland|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C379|ThymusGland|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C379|ThymusGland|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C379|ThymusGland|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C379|ThymusGland|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C379|ThymusGland|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C379|ThymusGland|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C379|ThymusGland|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C379|ThymusGland|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C379|ThymusGland|858|MalignantThymoma|8580/3|MalignantThymoma
C379|ThymusGland|858|MalignantThymoma|8581/3|MalignantTypeAThymoma
C379|ThymusGland|858|MalignantThymoma|8582/3|MalignantTypeABThymoma
C379|ThymusGland|858|MalignantThymoma|8583/3|MalignantTypeB1Thymoma
C379|ThymusGland|858|MalignantThymoma|8584/3|MalignantTypeB2Thymoma
C379|ThymusGland|858|MalignantThymoma|8585/3|ThymomaTypeB3
C379|ThymusGland|858|MalignantThymoma|8586/3|ThymicCarcinoma
C379|ThymusGland|858|MalignantThymoma|8588/3|NeoplasticEpithelialSpindleCell
C379|ThymusGland|858|MalignantThymoma|8589/3|CarcinomaShowingThymuslikeElement
C379|ThymusGland|908|Teratoma|9086/3|HematopoieticNeoplasm
C379|ThymusGland|959|Lymphoma|9590/3|Lymphoma
C379|ThymusGland|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C379|ThymusGland|959|Lymphoma|9596/3|CompositeLymphoma
C379|ThymusGland|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C379|ThymusGland|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C379|ThymusGland|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C379|ThymusGland|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C379|ThymusGland|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C379|ThymusGland|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C379|ThymusGland|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C379|ThymusGland|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C379|ThymusGland|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C379|ThymusGland|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C379|ThymusGland|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C379|ThymusGland|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C379|ThymusGland|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C379|ThymusGland|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C379|ThymusGland|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C379|ThymusGland|967|BCellLymphomas|9673/3|MantleCellLymphoma
C379|ThymusGland|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C379|ThymusGland|967|BCellLymphomas|9679/3|MediastinalLargeBcellLymphoma
C379|ThymusGland|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C379|ThymusGland|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C379|ThymusGland|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C379|ThymusGland|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C379|ThymusGland|969|FollicularAdenoma|9690/3|LymphomaFollicular
C379|ThymusGland|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C379|ThymusGland|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C379|ThymusGland|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C379|ThymusGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C379|ThymusGland|970|TCellLymphoma|9701/3|SezarySyndrome
C379|ThymusGland|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C379|ThymusGland|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C379|ThymusGland|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C379|ThymusGland|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C379|ThymusGland|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C379|ThymusGland|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C379|ThymusGland|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C379|ThymusGland|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C379|ThymusGland|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C379|ThymusGland|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C379|ThymusGland|973|Plasmacytoma|9731/3|Plasmacytoma
C379|ThymusGland|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C379|ThymusGland|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C379|ThymusGland|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C379|ThymusGland|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C379|ThymusGland|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C379|ThymusGland|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C379|ThymusGland|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C379|ThymusGland|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C379|ThymusGland|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C379|ThymusGland|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C379|ThymusGland|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C379|ThymusGland|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C379|ThymusGland|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C379|ThymusGland|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C379|ThymusGland|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C379|ThymusGland|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9812/3|null
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9813/3|null
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9814/3|null
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9817/3|null
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9818/3|null
C379|ThymusGland|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C379|ThymusGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C379|ThymusGland|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C379|ThymusGland|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C379|ThymusGland|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C379|ThymusGland|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C379|ThymusGland|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C379|ThymusGland|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C380|Heart|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C380|Heart|913|Hemangioendothelioma|9137/3|IntimalSarcoma
C380|Heart|959|Lymphoma|9590/3|Lymphoma
C380|Heart|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C380|Heart|959|Lymphoma|9596/3|CompositeLymphoma
C380|Heart|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C380|Heart|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C380|Heart|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C380|Heart|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C380|Heart|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C380|Heart|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C380|Heart|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C380|Heart|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C380|Heart|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C380|Heart|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C380|Heart|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C380|Heart|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C380|Heart|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C380|Heart|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C380|Heart|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C380|Heart|967|BCellLymphomas|9673/3|MantleCellLymphoma
C380|Heart|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C380|Heart|967|BCellLymphomas|9678/3|PrimaryEffusionLymphoma
C380|Heart|967|BCellLymphomas|9679/3|MediastinalLargeBcellLymphoma
C380|Heart|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C380|Heart|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C380|Heart|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C380|Heart|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C380|Heart|968|DiffuseLargeBCellLymphoma|9689/3|MucosaassociatedLymphoma
C380|Heart|969|FollicularAdenoma|9690/3|LymphomaFollicular
C380|Heart|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C380|Heart|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C380|Heart|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C380|Heart|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C380|Heart|970|TCellLymphoma|9700/3|MycosisFungoides
C380|Heart|970|TCellLymphoma|9701/3|SezarySyndrome
C380|Heart|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C380|Heart|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C380|Heart|970|TCellLymphoma|9708/3|TCellLymphoma
C380|Heart|970|TCellLymphoma|9709/3|CutaneousTCellNonHodgkinLymphoma
C380|Heart|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C380|Heart|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C380|Heart|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C380|Heart|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C380|Heart|971|AdultNonHodgkinLymphoma|9717/3|IntestinalTCellLymphomaNOS
C380|Heart|971|AdultNonHodgkinLymphoma|9718/3|CALCL
C380|Heart|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C380|Heart|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C380|Heart|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C380|Heart|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C380|Heart|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C380|Heart|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C380|Heart|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C380|Heart|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C380|Heart|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C380|Heart|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C380|Heart|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C380|Heart|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C380|Heart|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C380|Heart|981|PrecursorLymphoidNeoplasm|9812/3|null
C380|Heart|981|PrecursorLymphoidNeoplasm|9813/3|null
C380|Heart|981|PrecursorLymphoidNeoplasm|9814/3|null
C380|Heart|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C380|Heart|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C380|Heart|981|PrecursorLymphoidNeoplasm|9817/3|null
C380|Heart|981|PrecursorLymphoidNeoplasm|9818/3|null
C380|Heart|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C380|Heart|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C380|Heart|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C380|Heart|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C380|Heart|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C380|Heart|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C380|Heart|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C380|Heart|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C381-C383, C388|Mediastinum|868|Paraganglioma|8680/3|MalignantParaganglioma
C381-C383, C388|Mediastinum|869|MalignantExtraAdrenalParaganglioma|8693/3|MalignantExtraAdrenalParaganglioma
C381-C383, C388|Mediastinum|880|Sarcoma|8800/3|Sarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8801/3|SpindleCellSarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8802/3|GiantCellSarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8803/3|SmallCellSarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8804/3|SarcomaEpithelioid
C381-C383, C388|Mediastinum|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C381-C383, C388|Mediastinum|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C381-C383, C388|Mediastinum|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C381-C383, C388|Mediastinum|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C381-C383, C388|Mediastinum|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C381-C383, C388|Mediastinum|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C381-C383, C388|Mediastinum|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C381-C383, C388|Mediastinum|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8850/3|Liposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C381-C383, C388|Mediastinum|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8855/3|Liposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C381-C383, C388|Mediastinum|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C381-C383, C388|Mediastinum|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C381-C383, C388|Mediastinum|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C381-C383, C388|Mediastinum|889|MyomatousNeoplasm|8895/3|Myosarcoma
C381-C383, C388|Mediastinum|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C381-C383, C388|Mediastinum|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C381-C383, C388|Mediastinum|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C381-C383, C388|Mediastinum|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C381-C383, C388|Mediastinum|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C381-C383, C388|Mediastinum|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C381-C383, C388|Mediastinum|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C381-C383, C388|Mediastinum|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C381-C383, C388|Mediastinum|906|GermCellTumor|9060/3|Dysgerminoma
C381-C383, C388|Mediastinum|906|GermCellTumor|9061/3|Seminoma
C381-C383, C388|Mediastinum|906|GermCellTumor|9062/3|AtypicalSeminoma
C381-C383, C388|Mediastinum|906|GermCellTumor|9063/3|TesticularSpermatocyticSeminoma
C381-C383, C388|Mediastinum|906|GermCellTumor|9064/3|Germinoma
C381-C383, C388|Mediastinum|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C381-C383, C388|Mediastinum|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C381-C383, C388|Mediastinum|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C381-C383, C388|Mediastinum|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C381-C383, C388|Mediastinum|908|Teratoma|9080/3|ImmatureTeratoma
C381-C383, C388|Mediastinum|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C381-C383, C388|Mediastinum|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C381-C383, C388|Mediastinum|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C381-C383, C388|Mediastinum|908|Teratoma|9084/3|Teratoma
C381-C383, C388|Mediastinum|908|Teratoma|9085/3|MixedGermCellTumor
C381-C383, C388|Mediastinum|910|Choriocarcinoma|9100/3|Choriocarcinoma
C381-C383, C388|Mediastinum|910|Choriocarcinoma|9101/3|Choriocarcinoma
C381-C383, C388|Mediastinum|910|Choriocarcinoma|9105/3|EpithelioidTrophoblasticTumor
C381-C383, C388|Mediastinum|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9500/3|Neuroblastoma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9501/3|Medulloepithelioma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9503/3|Neuroepithelioma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C381-C383, C388|Mediastinum|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C381-C383, C388|Mediastinum|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C381-C383, C388|Mediastinum|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C381-C383, C388|Mediastinum|957|Perineurioma|9571/3|MalignantPerineurioma
C381-C383, C388|Mediastinum|959|Lymphoma|9590/3|Lymphoma
C381-C383, C388|Mediastinum|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C381-C383, C388|Mediastinum|959|Lymphoma|9596/3|CompositeLymphoma
C381-C383, C388|Mediastinum|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C381-C383, C388|Mediastinum|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C381-C383, C388|Mediastinum|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C381-C383, C388|Mediastinum|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C381-C383, C388|Mediastinum|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C381-C383, C388|Mediastinum|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C381-C383, C388|Mediastinum|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C381-C383, C388|Mediastinum|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C381-C383, C388|Mediastinum|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C381-C383, C388|Mediastinum|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C381-C383, C388|Mediastinum|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C381-C383, C388|Mediastinum|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C381-C383, C388|Mediastinum|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C381-C383, C388|Mediastinum|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C381-C383, C388|Mediastinum|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C381-C383, C388|Mediastinum|967|BCellLymphomas|9673/3|MantleCellLymphoma
C381-C383, C388|Mediastinum|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C381-C383, C388|Mediastinum|967|BCellLymphomas|9678/3|PrimaryEffusionLymphoma
C381-C383, C388|Mediastinum|967|BCellLymphomas|9679/3|MediastinalLargeBcellLymphoma
C381-C383, C388|Mediastinum|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C381-C383, C388|Mediastinum|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C381-C383, C388|Mediastinum|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C381-C383, C388|Mediastinum|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C381-C383, C388|Mediastinum|969|FollicularAdenoma|9690/3|LymphomaFollicular
C381-C383, C388|Mediastinum|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C381-C383, C388|Mediastinum|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C381-C383, C388|Mediastinum|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C381-C383, C388|Mediastinum|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C381-C383, C388|Mediastinum|970|TCellLymphoma|9701/3|SezarySyndrome
C381-C383, C388|Mediastinum|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C381-C383, C388|Mediastinum|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C381-C383, C388|Mediastinum|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C381-C383, C388|Mediastinum|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C381-C383, C388|Mediastinum|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C381-C383, C388|Mediastinum|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C381-C383, C388|Mediastinum|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C381-C383, C388|Mediastinum|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C381-C383, C388|Mediastinum|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C381-C383, C388|Mediastinum|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C381-C383, C388|Mediastinum|973|Plasmacytoma|9731/3|Plasmacytoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C381-C383, C388|Mediastinum|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C381-C383, C388|Mediastinum|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C381-C383, C388|Mediastinum|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C381-C383, C388|Mediastinum|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C381-C383, C388|Mediastinum|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C381-C383, C388|Mediastinum|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C381-C383, C388|Mediastinum|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C381-C383, C388|Mediastinum|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C381-C383, C388|Mediastinum|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C381-C383, C388|Mediastinum|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C381-C383, C388|Mediastinum|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C381-C383, C388|Mediastinum|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9812/3|null
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9813/3|null
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9814/3|null
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9817/3|null
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9818/3|null
C381-C383, C388|Mediastinum|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C381-C383, C388|Mediastinum|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C381-C383, C388|Mediastinum|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C381-C383, C388|Mediastinum|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C381-C383, C388|Mediastinum|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C381-C383, C388|Mediastinum|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C381-C383, C388|Mediastinum|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C381-C383, C388|Mediastinum|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C384|Pleura|880|Sarcoma|8800/3|Sarcoma
C384|Pleura|880|Sarcoma|8801/3|SpindleCellSarcoma
C384|Pleura|880|Sarcoma|8802/3|GiantCellSarcoma
C384|Pleura|880|Sarcoma|8803/3|SmallCellSarcoma
C384|Pleura|880|Sarcoma|8804/3|SarcomaEpithelioid
C384|Pleura|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C384|Pleura|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C384|Pleura|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C384|Pleura|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C384|Pleura|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C384|Pleura|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C384|Pleura|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C384|Pleura|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C384|Pleura|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C384|Pleura|897|Hepatoblastoma|8973/3|PleuropulmonaryBlastoma
C384|Pleura|905|MalignantMesothelioma|9050/3|MalignantMesothelioma
C384|Pleura|905|MalignantMesothelioma|9051/3|SarcomatoidMesothelioma
C384|Pleura|905|MalignantMesothelioma|9052/3|Mesothelioma
C384|Pleura|905|MalignantMesothelioma|9053/3|BiphasicMesothelioma
C384|Pleura|959|Lymphoma|9590/3|Lymphoma
C384|Pleura|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C384|Pleura|959|Lymphoma|9596/3|CompositeLymphoma
C384|Pleura|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C384|Pleura|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C384|Pleura|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C384|Pleura|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C384|Pleura|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C384|Pleura|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C384|Pleura|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C384|Pleura|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C384|Pleura|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C384|Pleura|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C384|Pleura|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C384|Pleura|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C384|Pleura|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C384|Pleura|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C384|Pleura|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C384|Pleura|967|BCellLymphomas|9673/3|MantleCellLymphoma
C384|Pleura|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C384|Pleura|967|BCellLymphomas|9678/3|PrimaryEffusionLymphoma
C384|Pleura|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C384|Pleura|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C384|Pleura|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C384|Pleura|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C384|Pleura|969|FollicularAdenoma|9690/3|LymphomaFollicular
C384|Pleura|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C384|Pleura|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C384|Pleura|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C384|Pleura|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C384|Pleura|970|TCellLymphoma|9701/3|SezarySyndrome
C384|Pleura|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C384|Pleura|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C384|Pleura|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C384|Pleura|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C384|Pleura|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C384|Pleura|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C384|Pleura|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C384|Pleura|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C384|Pleura|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C384|Pleura|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C384|Pleura|973|Plasmacytoma|9731/3|Plasmacytoma
C384|Pleura|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C384|Pleura|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C384|Pleura|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C384|Pleura|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C384|Pleura|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C384|Pleura|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C384|Pleura|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C384|Pleura|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C384|Pleura|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C384|Pleura|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C384|Pleura|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C384|Pleura|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C384|Pleura|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C384|Pleura|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C384|Pleura|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C384|Pleura|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C384|Pleura|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C384|Pleura|981|PrecursorLymphoidNeoplasm|9812/3|null
C384|Pleura|981|PrecursorLymphoidNeoplasm|9813/3|null
C384|Pleura|981|PrecursorLymphoidNeoplasm|9814/3|null
C384|Pleura|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C384|Pleura|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C384|Pleura|981|PrecursorLymphoidNeoplasm|9817/3|null
C384|Pleura|981|PrecursorLymphoidNeoplasm|9818/3|null
C384|Pleura|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C384|Pleura|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C384|Pleura|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C384|Pleura|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C384|Pleura|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C384|Pleura|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C384|Pleura|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C384|Pleura|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C390,C398-C399|RespiratorySystem|801|Carcinoma|8010/2|InSituCancer
C390,C398-C399|RespiratorySystem|801|Carcinoma|8010/3|CarcinomaNOSDNE
C390,C398-C399|RespiratorySystem|801|Carcinoma|8011/3|MalignantEpithelioma
C390,C398-C399|RespiratorySystem|801|Carcinoma|8012/3|LargeCellCarcinoma
C390,C398-C399|RespiratorySystem|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C390,C398-C399|RespiratorySystem|801|Carcinoma|8014/3|LargeCellCarcinoma
C390,C398-C399|RespiratorySystem|801|Carcinoma|8015/3|GlassyCellCarcinoma
C390,C398-C399|RespiratorySystem|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C390,C398-C399|RespiratorySystem|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C390,C398-C399|RespiratorySystem|802|Carcinoma|8022/3|PleomorphicCarcinoma
C390,C398-C399|RespiratorySystem|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C390,C398-C399|RespiratorySystem|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C390,C398-C399|RespiratorySystem|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C390,C398-C399|RespiratorySystem|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C390,C398-C399|RespiratorySystem|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C390,C398-C399|RespiratorySystem|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C390,C398-C399|RespiratorySystem|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C390,C398-C399|RespiratorySystem|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C390,C398-C399|RespiratorySystem|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C390,C398-C399|RespiratorySystem|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C390,C398-C399|RespiratorySystem|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C390,C398-C399|RespiratorySystem|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C390,C398-C399|RespiratorySystem|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C390,C398-C399|RespiratorySystem|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C390,C398-C399|RespiratorySystem|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C390,C398-C399|RespiratorySystem|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C390,C398-C399|RespiratorySystem|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C390,C398-C399|RespiratorySystem|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C390,C398-C399|RespiratorySystem|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C390,C398-C399|RespiratorySystem|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C390,C398-C399|RespiratorySystem|814|Adenocarcinoma|8140/3|Adenocarcinoma
C390,C398-C399|RespiratorySystem|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C390,C398-C399|RespiratorySystem|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C390,C398-C399|RespiratorySystem|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C390,C398-C399|RespiratorySystem|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C390,C398-C399|RespiratorySystem|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C390,C398-C399|RespiratorySystem|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C390,C398-C399|RespiratorySystem|823|SolidCarcinoma|8230/2|InSituCancer
C390,C398-C399|RespiratorySystem|823|SolidCarcinoma|8230/3|SolidCarcinoma
C390,C398-C399|RespiratorySystem|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C390,C398-C399|RespiratorySystem|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C390,C398-C399|RespiratorySystem|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C390,C398-C399|RespiratorySystem|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C390,C398-C399|RespiratorySystem|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C390,C398-C399|RespiratorySystem|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C390,C398-C399|RespiratorySystem|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C390,C398-C399|RespiratorySystem|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C390,C398-C399|RespiratorySystem|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C390,C398-C399|RespiratorySystem|825|BronchioloalveolarAdenocarcinoma|8250/3|LepidicPredominantAdenocarcinoma
C390,C398-C399|RespiratorySystem|825|BronchioloalveolarAdenocarcinoma|8251/3|BronchioloalveolarAdenocarcinoma
C390,C398-C399|RespiratorySystem|825|BronchioloalveolarAdenocarcinoma|8252/3|NonMucinousLungAdenocarcinomaInSitu
C390,C398-C399|RespiratorySystem|825|BronchioloalveolarAdenocarcinoma|8253/3|MucinousAdenocarcinoma
C390,C398-C399|RespiratorySystem|825|BronchioloalveolarAdenocarcinoma|8254/3|MixedSubtypeAdenocarcinomaOfLung
C390,C398-C399|RespiratorySystem|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C390,C398-C399|RespiratorySystem|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C390,C398-C399|RespiratorySystem|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C390,C398-C399|RespiratorySystem|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C390,C398-C399|RespiratorySystem|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C390,C398-C399|RespiratorySystem|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C390,C398-C399|RespiratorySystem|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C390,C398-C399|RespiratorySystem|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C390,C398-C399|RespiratorySystem|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C390,C398-C399|RespiratorySystem|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C390,C398-C399|RespiratorySystem|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C390,C398-C399|RespiratorySystem|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C390,C398-C399|RespiratorySystem|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C390,C398-C399|RespiratorySystem|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C390,C398-C399|RespiratorySystem|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C390,C398-C399|RespiratorySystem|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C390,C398-C399|RespiratorySystem|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C390,C398-C399|RespiratorySystem|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C390,C398-C399|RespiratorySystem|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C390,C398-C399|RespiratorySystem|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C390,C398-C399|RespiratorySystem|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C390,C398-C399|RespiratorySystem|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C390,C398-C399|RespiratorySystem|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C390,C398-C399|RespiratorySystem|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C390,C398-C399|RespiratorySystem|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C390,C398-C399|RespiratorySystem|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C390,C398-C399|RespiratorySystem|880|Sarcoma|8800/3|Sarcoma
C390,C398-C399|RespiratorySystem|880|Sarcoma|8801/3|SpindleCellSarcoma
C390,C398-C399|RespiratorySystem|880|Sarcoma|8802/3|GiantCellSarcoma
C390,C398-C399|RespiratorySystem|880|Sarcoma|8803/3|SmallCellSarcoma
C390,C398-C399|RespiratorySystem|880|Sarcoma|8804/3|SarcomaEpithelioid
C390,C398-C399|RespiratorySystem|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C390,C398-C399|RespiratorySystem|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C390,C398-C399|RespiratorySystem|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C390,C398-C399|RespiratorySystem|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C390,C398-C399|RespiratorySystem|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C390,C398-C399|RespiratorySystem|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C390,C398-C399|RespiratorySystem|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C390,C398-C399|RespiratorySystem|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C390,C398-C399|RespiratorySystem|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C390,C398-C399|RespiratorySystem|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C390,C398-C399|RespiratorySystem|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C390,C398-C399|RespiratorySystem|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C390,C398-C399|RespiratorySystem|889|MyomatousNeoplasm|8895/3|Myosarcoma
C390,C398-C399|RespiratorySystem|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C390,C398-C399|RespiratorySystem|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C390,C398-C399|RespiratorySystem|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C390,C398-C399|RespiratorySystem|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C390,C398-C399|RespiratorySystem|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C390,C398-C399|RespiratorySystem|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C390,C398-C399|RespiratorySystem|898|Carcinosarcoma|8980/3|Carcinosarcoma
C390,C398-C399|RespiratorySystem|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C390,C398-C399|RespiratorySystem|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C390,C398-C399|RespiratorySystem|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C390,C398-C399|RespiratorySystem|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C390,C398-C399|RespiratorySystem|908|Teratoma|9080/3|ImmatureTeratoma
C390,C398-C399|RespiratorySystem|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C390,C398-C399|RespiratorySystem|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C390,C398-C399|RespiratorySystem|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C390,C398-C399|RespiratorySystem|908|Teratoma|9084/3|Teratoma
C390,C398-C399|RespiratorySystem|908|Teratoma|9085/3|MixedGermCellTumor
C390,C398-C399|RespiratorySystem|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C390,C398-C399|RespiratorySystem|936|NeuroepitheliomaPeripheral|9364/3|NeuroepitheliomaPeripheral
C390,C398-C399|RespiratorySystem|936|NeuroepitheliomaPeripheral|9365/3|AskinTumor
C390,C398-C399|RespiratorySystem|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8800/3|Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8801/3|SpindleCellSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8802/3|GiantCellSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8803/3|SmallCellSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8804/3|SarcomaEpithelioid
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|FibromatousNeoplasm|8812/3|PeriostealFibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|884|Myxosarcoma|8840/3|Myxosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8850/3|Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8855/3|Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|904|SynovialSarcoma|9040/3|SynovialSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|904|SynovialSarcoma|9041/3|SpindleCellSynovialSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|904|SynovialSarcoma|9042/3|EpithelialSynovialSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|904|SynovialSarcoma|9043/3|BiphasicSynovialSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9180/3|Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9181/3|ChondroblasticOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9182/3|FibroblasticOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9183/3|TelangiectaticOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9184/3|PagetDisease
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9185/3|SmallCellOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9186/3|ConventionalOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9187/3|Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|919|ParostealOsteosarcoma|9192/3|ParostealOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|919|ParostealOsteosarcoma|9193/3|PeriostealOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|919|ParostealOsteosarcoma|9194/3|HighGradeSurfaceOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|919|ParostealOsteosarcoma|9195/3|ConventionalOsteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|922|Chondrosarcoma|9220/3|Chondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|922|Chondrosarcoma|9221/3|PeriostealChondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|923|ChondroblastomaMalignant|9230/3|ChondroblastomaMalignant
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|923|ChondroblastomaMalignant|9231/3|MyxoidChondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|924|OsseousAndChondromatousNeoplasms|9240/3|MesenchymalChondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|924|OsseousAndChondromatousNeoplasms|9242/3|ClearCellChondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|924|OsseousAndChondromatousNeoplasms|9243/3|DedifferentiatedChondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|925|BoneNeoplasm|9250/3|GiantCellTumorOfBone
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|925|BoneNeoplasm|9251/3|GiantCellTumorOfSoftTissue
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|926|EwingSarcoma|9260/3|EwingSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|926|EwingSarcoma|9261/3|Adamantinoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|927|OdontogenicNeoplasm|9270/3|MalignantOdontogenicTumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|929|AmeloblasticOdontosarcoma|9290/3|AmeloblasticOdontosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|931|MalignantAmeloblastoma|9310/3|MalignantAmeloblastoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|933|AmeloblasticFibrosarcoma|9330/3|AmeloblasticFibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|934|MalignantOdontogenicTumor|9342/3|MalignantOdontogenicTumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|936|NeuroepitheliomaPeripheral|9364/3|NeuroepitheliomaPeripheral
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|936|NeuroepitheliomaPeripheral|9365/3|AskinTumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|937|Chordoma|9370/3|Chordoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|937|Chordoma|9371/3|ChondroidChordoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|937|Chordoma|9372/3|DedifferentiatedChordoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|959|Lymphoma|9590/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|959|Lymphoma|9596/3|CompositeLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|967|BCellLymphomas|9673/3|MantleCellLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|FollicularAdenoma|9690/3|LymphomaFollicular
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|970|TCellLymphoma|9701/3|SezarySyndrome
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9731/3|Plasmacytoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9732/3|PlasmaCellMyeloma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9812/3|null
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9813/3|null
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9814/3|null
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9817/3|null
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9818/3|null
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C410|Skull|880|Sarcoma|8800/3|Sarcoma
C410|Skull|880|Sarcoma|8801/3|SpindleCellSarcoma
C410|Skull|880|Sarcoma|8802/3|GiantCellSarcoma
C410|Skull|880|Sarcoma|8803/3|SmallCellSarcoma
C410|Skull|880|Sarcoma|8804/3|SarcomaEpithelioid
C410|Skull|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C410|Skull|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C410|Skull|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C410|Skull|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C410|Skull|881|FibromatousNeoplasm|8812/3|PeriostealFibrosarcoma
C410|Skull|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C410|Skull|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C410|Skull|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C410|Skull|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C410|Skull|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C410|Skull|884|Myxosarcoma|8840/3|Myxosarcoma
C410|Skull|885|Liposarcoma|8850/3|Liposarcoma
C410|Skull|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C410|Skull|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C410|Skull|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C410|Skull|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C410|Skull|885|Liposarcoma|8855/3|Liposarcoma
C410|Skull|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C410|Skull|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C410|Skull|904|SynovialSarcoma|9040/3|SynovialSarcoma
C410|Skull|904|SynovialSarcoma|9041/3|SpindleCellSynovialSarcoma
C410|Skull|904|SynovialSarcoma|9042/3|EpithelialSynovialSarcoma
C410|Skull|904|SynovialSarcoma|9043/3|BiphasicSynovialSarcoma
C410|Skull|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C410|Skull|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C410|Skull|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C410|Skull|918|Osteosarcoma|9180/3|Osteosarcoma
C410|Skull|918|Osteosarcoma|9181/3|ChondroblasticOsteosarcoma
C410|Skull|918|Osteosarcoma|9182/3|FibroblasticOsteosarcoma
C410|Skull|918|Osteosarcoma|9183/3|TelangiectaticOsteosarcoma
C410|Skull|918|Osteosarcoma|9184/3|PagetDisease
C410|Skull|918|Osteosarcoma|9185/3|SmallCellOsteosarcoma
C410|Skull|918|Osteosarcoma|9186/3|ConventionalOsteosarcoma
C410|Skull|918|Osteosarcoma|9187/3|Osteosarcoma
C410|Skull|919|ParostealOsteosarcoma|9192/3|ParostealOsteosarcoma
C410|Skull|919|ParostealOsteosarcoma|9193/3|PeriostealOsteosarcoma
C410|Skull|919|ParostealOsteosarcoma|9194/3|HighGradeSurfaceOsteosarcoma
C410|Skull|919|ParostealOsteosarcoma|9195/3|ConventionalOsteosarcoma
C410|Skull|922|Chondrosarcoma|9220/3|Chondrosarcoma
C410|Skull|922|Chondrosarcoma|9221/3|PeriostealChondrosarcoma
C410|Skull|923|ChondroblastomaMalignant|9230/3|ChondroblastomaMalignant
C410|Skull|923|ChondroblastomaMalignant|9231/3|MyxoidChondrosarcoma
C410|Skull|924|OsseousAndChondromatousNeoplasms|9240/3|MesenchymalChondrosarcoma
C410|Skull|924|OsseousAndChondromatousNeoplasms|9242/3|ClearCellChondrosarcoma
C410|Skull|924|OsseousAndChondromatousNeoplasms|9243/3|DedifferentiatedChondrosarcoma
C410|Skull|925|BoneNeoplasm|9250/3|GiantCellTumorOfBone
C410|Skull|925|BoneNeoplasm|9251/3|GiantCellTumorOfSoftTissue
C410|Skull|926|EwingSarcoma|9260/3|EwingSarcoma
C410|Skull|926|EwingSarcoma|9261/3|Adamantinoma
C410|Skull|927|OdontogenicNeoplasm|9270/3|MalignantOdontogenicTumor
C410|Skull|929|AmeloblasticOdontosarcoma|9290/3|AmeloblasticOdontosarcoma
C410|Skull|930|OdontogenicNeoplasm|9302/3|GhostCellOdontogenicCarcinoma
C410|Skull|931|MalignantAmeloblastoma|9310/3|MalignantAmeloblastoma
C410|Skull|933|AmeloblasticFibrosarcoma|9330/3|AmeloblasticFibrosarcoma
C410|Skull|934|MalignantOdontogenicTumor|9341/3|ClearCellOdontogenicCarcinoma
C410|Skull|934|MalignantOdontogenicTumor|9342/3|MalignantOdontogenicTumor
C410|Skull|936|NeuroepitheliomaPeripheral|9364/3|NeuroepitheliomaPeripheral
C410|Skull|936|NeuroepitheliomaPeripheral|9365/3|AskinTumor
C410|Skull|937|Chordoma|9370/3|Chordoma
C410|Skull|937|Chordoma|9371/3|ChondroidChordoma
C410|Skull|937|Chordoma|9372/3|DedifferentiatedChordoma
C410|Skull|959|Lymphoma|9590/3|Lymphoma
C410|Skull|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C410|Skull|959|Lymphoma|9596/3|CompositeLymphoma
C410|Skull|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C410|Skull|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C410|Skull|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C410|Skull|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C410|Skull|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C410|Skull|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C410|Skull|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C410|Skull|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C410|Skull|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C410|Skull|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C410|Skull|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C410|Skull|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C410|Skull|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C410|Skull|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C410|Skull|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C410|Skull|967|BCellLymphomas|9673/3|MantleCellLymphoma
C410|Skull|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C410|Skull|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C410|Skull|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C410|Skull|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C410|Skull|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C410|Skull|969|FollicularAdenoma|9690/3|LymphomaFollicular
C410|Skull|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C410|Skull|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C410|Skull|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C410|Skull|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C410|Skull|970|TCellLymphoma|9701/3|SezarySyndrome
C410|Skull|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C410|Skull|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C410|Skull|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C410|Skull|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C410|Skull|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C410|Skull|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C410|Skull|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C410|Skull|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C410|Skull|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C410|Skull|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C410|Skull|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C410|Skull|973|Plasmacytoma|9731/3|Plasmacytoma
C410|Skull|973|Plasmacytoma|9732/3|PlasmaCellMyeloma
C410|Skull|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C410|Skull|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C410|Skull|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C410|Skull|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C410|Skull|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C410|Skull|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C410|Skull|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C410|Skull|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C410|Skull|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C410|Skull|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C410|Skull|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C410|Skull|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C410|Skull|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C410|Skull|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C410|Skull|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C410|Skull|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C410|Skull|981|PrecursorLymphoidNeoplasm|9812/3|null
C410|Skull|981|PrecursorLymphoidNeoplasm|9813/3|null
C410|Skull|981|PrecursorLymphoidNeoplasm|9814/3|null
C410|Skull|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C410|Skull|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C410|Skull|981|PrecursorLymphoidNeoplasm|9817/3|null
C410|Skull|981|PrecursorLymphoidNeoplasm|9818/3|null
C410|Skull|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C410|Skull|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C410|Skull|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C410|Skull|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C410|Skull|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C410|Skull|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C410|Skull|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C410|Skull|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C411|Mandible|880|Sarcoma|8800/3|Sarcoma
C411|Mandible|880|Sarcoma|8801/3|SpindleCellSarcoma
C411|Mandible|880|Sarcoma|8802/3|GiantCellSarcoma
C411|Mandible|880|Sarcoma|8803/3|SmallCellSarcoma
C411|Mandible|880|Sarcoma|8804/3|SarcomaEpithelioid
C411|Mandible|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C411|Mandible|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C411|Mandible|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C411|Mandible|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C411|Mandible|881|FibromatousNeoplasm|8812/3|PeriostealFibrosarcoma
C411|Mandible|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C411|Mandible|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C411|Mandible|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C411|Mandible|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C411|Mandible|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C411|Mandible|884|Myxosarcoma|8840/3|Myxosarcoma
C411|Mandible|885|Liposarcoma|8850/3|Liposarcoma
C411|Mandible|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C411|Mandible|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C411|Mandible|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C411|Mandible|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C411|Mandible|885|Liposarcoma|8855/3|Liposarcoma
C411|Mandible|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C411|Mandible|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C411|Mandible|904|SynovialSarcoma|9040/3|SynovialSarcoma
C411|Mandible|904|SynovialSarcoma|9041/3|SpindleCellSynovialSarcoma
C411|Mandible|904|SynovialSarcoma|9042/3|EpithelialSynovialSarcoma
C411|Mandible|904|SynovialSarcoma|9043/3|BiphasicSynovialSarcoma
C411|Mandible|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C411|Mandible|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C411|Mandible|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C411|Mandible|918|Osteosarcoma|9180/3|Osteosarcoma
C411|Mandible|918|Osteosarcoma|9181/3|ChondroblasticOsteosarcoma
C411|Mandible|918|Osteosarcoma|9182/3|FibroblasticOsteosarcoma
C411|Mandible|918|Osteosarcoma|9183/3|TelangiectaticOsteosarcoma
C411|Mandible|918|Osteosarcoma|9184/3|PagetDisease
C411|Mandible|918|Osteosarcoma|9185/3|SmallCellOsteosarcoma
C411|Mandible|918|Osteosarcoma|9186/3|ConventionalOsteosarcoma
C411|Mandible|918|Osteosarcoma|9187/3|Osteosarcoma
C411|Mandible|919|ParostealOsteosarcoma|9192/3|ParostealOsteosarcoma
C411|Mandible|919|ParostealOsteosarcoma|9193/3|PeriostealOsteosarcoma
C411|Mandible|919|ParostealOsteosarcoma|9194/3|HighGradeSurfaceOsteosarcoma
C411|Mandible|919|ParostealOsteosarcoma|9195/3|ConventionalOsteosarcoma
C411|Mandible|922|Chondrosarcoma|9220/3|Chondrosarcoma
C411|Mandible|922|Chondrosarcoma|9221/3|PeriostealChondrosarcoma
C411|Mandible|923|ChondroblastomaMalignant|9230/3|ChondroblastomaMalignant
C411|Mandible|923|ChondroblastomaMalignant|9231/3|MyxoidChondrosarcoma
C411|Mandible|924|OsseousAndChondromatousNeoplasms|9240/3|MesenchymalChondrosarcoma
C411|Mandible|924|OsseousAndChondromatousNeoplasms|9242/3|ClearCellChondrosarcoma
C411|Mandible|924|OsseousAndChondromatousNeoplasms|9243/3|DedifferentiatedChondrosarcoma
C411|Mandible|925|BoneNeoplasm|9250/3|GiantCellTumorOfBone
C411|Mandible|925|BoneNeoplasm|9251/3|GiantCellTumorOfSoftTissue
C411|Mandible|926|EwingSarcoma|9260/3|EwingSarcoma
C411|Mandible|926|EwingSarcoma|9261/3|Adamantinoma
C411|Mandible|927|OdontogenicNeoplasm|9270/3|MalignantOdontogenicTumor
C411|Mandible|929|AmeloblasticOdontosarcoma|9290/3|AmeloblasticOdontosarcoma
C411|Mandible|930|OdontogenicNeoplasm|9302/3|GhostCellOdontogenicCarcinoma
C411|Mandible|931|MalignantAmeloblastoma|9310/3|MalignantAmeloblastoma
C411|Mandible|933|AmeloblasticFibrosarcoma|9330/3|AmeloblasticFibrosarcoma
C411|Mandible|934|MalignantOdontogenicTumor|9341/3|ClearCellOdontogenicCarcinoma
C411|Mandible|934|MalignantOdontogenicTumor|9342/3|MalignantOdontogenicTumor
C411|Mandible|936|NeuroepitheliomaPeripheral|9364/3|NeuroepitheliomaPeripheral
C411|Mandible|936|NeuroepitheliomaPeripheral|9365/3|AskinTumor
C411|Mandible|937|Chordoma|9370/3|Chordoma
C411|Mandible|937|Chordoma|9371/3|ChondroidChordoma
C411|Mandible|937|Chordoma|9372/3|DedifferentiatedChordoma
C411|Mandible|959|Lymphoma|9590/3|Lymphoma
C411|Mandible|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C411|Mandible|959|Lymphoma|9596/3|CompositeLymphoma
C411|Mandible|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C411|Mandible|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C411|Mandible|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C411|Mandible|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C411|Mandible|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C411|Mandible|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C411|Mandible|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C411|Mandible|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C411|Mandible|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C411|Mandible|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C411|Mandible|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C411|Mandible|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C411|Mandible|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C411|Mandible|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C411|Mandible|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C411|Mandible|967|BCellLymphomas|9673/3|MantleCellLymphoma
C411|Mandible|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C411|Mandible|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C411|Mandible|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C411|Mandible|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C411|Mandible|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C411|Mandible|969|FollicularAdenoma|9690/3|LymphomaFollicular
C411|Mandible|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C411|Mandible|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C411|Mandible|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C411|Mandible|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C411|Mandible|970|TCellLymphoma|9701/3|SezarySyndrome
C411|Mandible|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C411|Mandible|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C411|Mandible|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C411|Mandible|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C411|Mandible|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C411|Mandible|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C411|Mandible|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C411|Mandible|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C411|Mandible|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C411|Mandible|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C411|Mandible|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C411|Mandible|973|Plasmacytoma|9731/3|Plasmacytoma
C411|Mandible|973|Plasmacytoma|9732/3|PlasmaCellMyeloma
C411|Mandible|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C411|Mandible|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C411|Mandible|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C411|Mandible|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C411|Mandible|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C411|Mandible|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C411|Mandible|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C411|Mandible|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C411|Mandible|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C411|Mandible|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C411|Mandible|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C411|Mandible|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C411|Mandible|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C411|Mandible|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C411|Mandible|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C411|Mandible|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C411|Mandible|981|PrecursorLymphoidNeoplasm|9812/3|null
C411|Mandible|981|PrecursorLymphoidNeoplasm|9813/3|null
C411|Mandible|981|PrecursorLymphoidNeoplasm|9814/3|null
C411|Mandible|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C411|Mandible|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C411|Mandible|981|PrecursorLymphoidNeoplasm|9817/3|null
C411|Mandible|981|PrecursorLymphoidNeoplasm|9818/3|null
C411|Mandible|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C411|Mandible|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C411|Mandible|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C411|Mandible|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C411|Mandible|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C411|Mandible|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C411|Mandible|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C411|Mandible|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C420, C421, C424|BoneMarrow|959|Lymphoma|9590/3|Lymphoma
C420, C421, C424|BoneMarrow|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C420, C421, C424|BoneMarrow|959|Lymphoma|9596/3|CompositeLymphoma
C420, C421, C424|BoneMarrow|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C420, C421, C424|BoneMarrow|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C420, C421, C424|BoneMarrow|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C420, C421, C424|BoneMarrow|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C420, C421, C424|BoneMarrow|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C420, C421, C424|BoneMarrow|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C420, C421, C424|BoneMarrow|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C420, C421, C424|BoneMarrow|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C420, C421, C424|BoneMarrow|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C420, C421, C424|BoneMarrow|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C420, C421, C424|BoneMarrow|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C420, C421, C424|BoneMarrow|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C420, C421, C424|BoneMarrow|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C420, C421, C424|BoneMarrow|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C420, C421, C424|BoneMarrow|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C420, C421, C424|BoneMarrow|967|BCellLymphomas|9673/3|MantleCellLymphoma
C420, C421, C424|BoneMarrow|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C420, C421, C424|BoneMarrow|967|BCellLymphomas|9678/3|PrimaryEffusionLymphoma
C420, C421, C424|BoneMarrow|967|BCellLymphomas|9679/3|MediastinalLargeBcellLymphoma
C420, C421, C424|BoneMarrow|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C420, C421, C424|BoneMarrow|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C420, C421, C424|BoneMarrow|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C420, C421, C424|BoneMarrow|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C420, C421, C424|BoneMarrow|968|DiffuseLargeBCellLymphoma|9689/3|MucosaassociatedLymphoma
C420, C421, C424|BoneMarrow|969|FollicularAdenoma|9690/3|LymphomaFollicular
C420, C421, C424|BoneMarrow|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C420, C421, C424|BoneMarrow|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C420, C421, C424|BoneMarrow|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C420, C421, C424|BoneMarrow|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C420, C421, C424|BoneMarrow|970|TCellLymphoma|9701/3|SezarySyndrome
C420, C421, C424|BoneMarrow|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C420, C421, C424|BoneMarrow|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C420, C421, C424|BoneMarrow|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C420, C421, C424|BoneMarrow|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C420, C421, C424|BoneMarrow|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C420, C421, C424|BoneMarrow|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C420, C421, C424|BoneMarrow|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C420, C421, C424|BoneMarrow|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C420, C421, C424|BoneMarrow|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C420, C421, C424|BoneMarrow|973|Plasmacytoma|9731/3|Plasmacytoma
C420, C421, C424|BoneMarrow|973|Plasmacytoma|9732/3|PlasmaCellMyeloma
C420, C421, C424|BoneMarrow|973|Plasmacytoma|9733/3|PlasmaCellLeukemia
C420, C421, C424|BoneMarrow|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C420, C421, C424|BoneMarrow|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C420, C421, C424|BoneMarrow|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C420, C421, C424|BoneMarrow|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C420, C421, C424|BoneMarrow|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C420, C421, C424|BoneMarrow|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C420, C421, C424|BoneMarrow|974|MastCellNeoplasm|9742/3|MastCellLeukemia
C420, C421, C424|BoneMarrow|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C420, C421, C424|BoneMarrow|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C420, C421, C424|BoneMarrow|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C420, C421, C424|BoneMarrow|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C420, C421, C424|BoneMarrow|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C420, C421, C424|BoneMarrow|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C420, C421, C424|BoneMarrow|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C420, C421, C424|BoneMarrow|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C420, C421, C424|BoneMarrow|976|ImmunoproliferativeDisorder|9760/3|ImmunoproliferativeDisorder
C420, C421, C424|BoneMarrow|976|ImmunoproliferativeDisorder|9761/3|WaldenstromMacroglobulinemia
C420, C421, C424|BoneMarrow|976|ImmunoproliferativeDisorder|9762/3|HeavyChainDisease
C420, C421, C424|BoneMarrow|980|Leukemia|9800/3|Leukemia
C420, C421, C424|BoneMarrow|980|Leukemia|9801/3|AcuteLeukemia
C420, C421, C424|BoneMarrow|980|Leukemia|9805/3|AcuteBiphenotypicLeukemia
C420, C421, C424|BoneMarrow|980|Leukemia|9806/3|MixedPhenotypeAcuteLeukemia
C420, C421, C424|BoneMarrow|980|Leukemia|9807/3|MixedPhenotypeAcuteLeukemia
C420, C421, C424|BoneMarrow|980|Leukemia|9808/3|MixedPhenotypeAcuteLeukemia
C420, C421, C424|BoneMarrow|980|Leukemia|9809/3|MixedPhenotypeAcuteLeukemia
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9812/3|null
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9813/3|null
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9814/3|null
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9817/3|null
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9818/3|null
C420, C421, C424|BoneMarrow|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C420, C421, C424|BoneMarrow|982|LymphoidLeukemia|9820/3|LymphoidLeukemia
C420, C421, C424|BoneMarrow|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C420, C421, C424|BoneMarrow|982|LymphoidLeukemia|9826/3|BurkittLeukemia
C420, C421, C424|BoneMarrow|982|LymphoidLeukemia|9827/3|AdultTcellLeukemia
C420, C421, C424|BoneMarrow|982|LymphoidLeukemia|9828/3|L2AcuteLymphoblasticLeukemia
C420, C421, C424|BoneMarrow|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C420, C421, C424|BoneMarrow|983|Leukemia|9832/3|ProlymphocyticLeukemia
C420, C421, C424|BoneMarrow|983|Leukemia|9833/3|BCellProlymphocyticLeukemia
C420, C421, C424|BoneMarrow|983|Leukemia|9834/3|TCellProlymphocyticLeukemia
C420, C421, C424|BoneMarrow|983|Leukemia|9835/3|AcuteLymphoblasticLeukemia
C420, C421, C424|BoneMarrow|983|Leukemia|9836/3|BAcuteLymphoblasticLeukemia
C420, C421, C424|BoneMarrow|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C420, C421, C424|BoneMarrow|984|Leukemia|9840/3|AcuteErythroidLeukemia
C420, C421, C424|BoneMarrow|986|MyeloidLeukemia|9860/3|MyeloidLeukemia
C420, C421, C424|BoneMarrow|986|MyeloidLeukemia|9861/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|986|MyeloidLeukemia|9863/3|MyeloidLeukemiaChronic
C420, C421, C424|BoneMarrow|986|MyeloidLeukemia|9865/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|986|MyeloidLeukemia|9866/3|AcutePromyelocyticLeukemia
C420, C421, C424|BoneMarrow|986|MyeloidLeukemia|9867/3|AcuteMyelomonocyticLeukemia
C420, C421, C424|BoneMarrow|986|MyeloidLeukemia|9869/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9870/3|AcuteBasophilicLeukemia
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9871/3|CMMLWithEosinophilia
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9872/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9873/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9874/3|AcuteMyeloidLeukemiaWithMaturation
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9875/3|MyeloidLeukemiaChronic
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9876/3|SubacuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9877/3|AcuteMyeloidLeukemiaWithMutatedNPM1
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9878/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|987|MyeloidLeukemia|9879/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|989|Leukemia|9891/3|AcuteMonocyticLeukemia
C420, C421, C424|BoneMarrow|989|Leukemia|9895/3|AMLWithMultilineageDysplasia
C420, C421, C424|BoneMarrow|989|Leukemia|9896/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|989|Leukemia|9897/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|989|Leukemia|9898/3|MyeloidLeukemia
C420, C421, C424|BoneMarrow|991|AcuteMegakaryocyticLeukemias|9910/3|AcuteMegakaryocyticLeukemias
C420, C421, C424|BoneMarrow|991|AcuteMegakaryocyticLeukemias|9911/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|991|AcuteMegakaryocyticLeukemias|9912/3|AcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|992|TherapyRelatedLeukemia|9920/3|TherapyRelatedAcuteMyeloidLeukemia
C420, C421, C424|BoneMarrow|993|MyeloidSarcoma|9930/3|MyeloidSarcoma
C420, C421, C424|BoneMarrow|993|MyeloidSarcoma|9931/3|AcutePanmyelosisWithMyelofibrosis
C420, C421, C424|BoneMarrow|994|Leukemia|9940/3|HairyCellLeukemia
C420, C421, C424|BoneMarrow|994|Leukemia|9945/3|ChronicMyelomonocyticLeukemia
C420, C421, C424|BoneMarrow|994|Leukemia|9946/3|JuvenileMyelomonocyticLeukemia
C420, C421, C424|BoneMarrow|994|Leukemia|9948/3|AggressiveNKCellLeukemia
C420, C421, C424|BoneMarrow|995|PolycythemiaVera|9950/3|PolycythemiaVera
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9960/3|MyeloproliferativeNeoplasm
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9961/3|PrimaryMyelofibrosis
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9962/3|EssentialThrombocythemia
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9963/3|ChronicNeutrophilicLeukemia
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9964/3|HypereosinophilicSyndrome
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9966/3|LymphocyticNeoplasm
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C420, C421, C424|BoneMarrow|996|MyeloproliferativeNeoplasm|9968/3|LymphocyticNeoplasm
C420, C421, C424|BoneMarrow|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C420, C421, C424|BoneMarrow|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C420, C421, C424|BoneMarrow|998|RefractoryAnemia|9980/3|RefractoryAnemia
C420, C421, C424|BoneMarrow|998|RefractoryAnemia|9982/3|RefractoryAnemiaWithSideroblasts
C420, C421, C424|BoneMarrow|998|RefractoryAnemia|9983/3|RefractoryAnemiaWithExcessBlasts
C420, C421, C424|BoneMarrow|998|RefractoryAnemia|9984/3|RefractoryAnemiaWithExcessBlasts
C420, C421, C424|BoneMarrow|998|RefractoryAnemia|9985/3|RefractoryCytopeniaOfChildhood
C420, C421, C424|BoneMarrow|998|RefractoryAnemia|9986/3|5qsyndrome
C420, C421, C424|BoneMarrow|998|RefractoryAnemia|9987/3|MyelodysplasticSyndrome
C420, C421, C424|BoneMarrow|998|RefractoryAnemia|9989/3|MyelodysplasticSyndrome
C420, C421, C424|BoneMarrow|999|MyelodysplasticSyndrome|9991/3|RefractoryNeutropenia
C420, C421, C424|BoneMarrow|999|MyelodysplasticSyndrome|9992/3|RefractoryThrombocytopenia
C420, C421, C424|BoneMarrow|999|MyelodysplasticSyndrome|9993/3|MyelodysplasticSyndrome
C422|Spleen|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C422|Spleen|959|Lymphoma|9590/3|Lymphoma
C422|Spleen|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C422|Spleen|959|Lymphoma|9596/3|CompositeLymphoma
C422|Spleen|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C422|Spleen|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C422|Spleen|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C422|Spleen|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C422|Spleen|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C422|Spleen|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C422|Spleen|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C422|Spleen|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C422|Spleen|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C422|Spleen|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C422|Spleen|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C422|Spleen|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C422|Spleen|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C422|Spleen|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C422|Spleen|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C422|Spleen|967|BCellLymphomas|9673/3|MantleCellLymphoma
C422|Spleen|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C422|Spleen|967|BCellLymphomas|9678/3|PrimaryEffusionLymphoma
C422|Spleen|967|BCellLymphomas|9679/3|MediastinalLargeBcellLymphoma
C422|Spleen|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C422|Spleen|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C422|Spleen|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C422|Spleen|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C422|Spleen|968|DiffuseLargeBCellLymphoma|9689/3|MucosaassociatedLymphoma
C422|Spleen|969|FollicularAdenoma|9690/3|LymphomaFollicular
C422|Spleen|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C422|Spleen|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C422|Spleen|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C422|Spleen|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C422|Spleen|970|TCellLymphoma|9701/3|SezarySyndrome
C422|Spleen|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C422|Spleen|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C422|Spleen|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C422|Spleen|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C422|Spleen|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C422|Spleen|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C422|Spleen|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C422|Spleen|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C422|Spleen|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C422|Spleen|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C422|Spleen|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C422|Spleen|973|Plasmacytoma|9731/3|Plasmacytoma
C422|Spleen|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C422|Spleen|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C422|Spleen|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C422|Spleen|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C422|Spleen|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C422|Spleen|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C422|Spleen|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C422|Spleen|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C422|Spleen|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C422|Spleen|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C422|Spleen|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C422|Spleen|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C422|Spleen|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C422|Spleen|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C422|Spleen|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C422|Spleen|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C422|Spleen|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C422|Spleen|981|PrecursorLymphoidNeoplasm|9812/3|null
C422|Spleen|981|PrecursorLymphoidNeoplasm|9813/3|null
C422|Spleen|981|PrecursorLymphoidNeoplasm|9814/3|null
C422|Spleen|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C422|Spleen|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C422|Spleen|981|PrecursorLymphoidNeoplasm|9817/3|null
C422|Spleen|981|PrecursorLymphoidNeoplasm|9818/3|null
C422|Spleen|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C422|Spleen|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C422|Spleen|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C422|Spleen|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C422|Spleen|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C422|Spleen|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C422|Spleen|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C422|Spleen|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C423|ReticuloendothelialSystem|959|Lymphoma|9590/3|Lymphoma
C423|ReticuloendothelialSystem|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C423|ReticuloendothelialSystem|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C423|ReticuloendothelialSystem|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C423|ReticuloendothelialSystem|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C423|ReticuloendothelialSystem|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C423|ReticuloendothelialSystem|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C423|ReticuloendothelialSystem|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C423|ReticuloendothelialSystem|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C423|ReticuloendothelialSystem|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C423|ReticuloendothelialSystem|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C440-C449|Skin|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C440-C449|Skin|811|PilomatricalCarcinoma|8110/3|PilomatricalCarcinoma
C440-C449|Skin|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C440-C449|Skin|814|Adenocarcinoma|8140/3|Adenocarcinoma
C440-C449|Skin|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C440-C449|Skin|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C440-C449|Skin|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C440-C449|Skin|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C440-C449|Skin|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C440-C449|Skin|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C440-C449|Skin|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C440-C449|Skin|823|SolidCarcinoma|8230/2|InSituCancer
C440-C449|Skin|823|SolidCarcinoma|8230/3|SolidCarcinoma
C440-C449|Skin|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C440-C449|Skin|824|AtypicalCarcinoidTumor|8247/3|MerkelCellCarcinoma
C440-C449|Skin|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C440-C449|Skin|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C440-C449|Skin|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C440-C449|Skin|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C440-C449|Skin|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C440-C449|Skin|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C440-C449|Skin|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C440-C449|Skin|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C440-C449|Skin|839|AdnexalCarcinoma|8390/3|AdnexalCarcinoma
C440-C449|Skin|840|SweatGlandAdenocarcinoma|8400/3|SweatGlandAdenocarcinoma
C440-C449|Skin|840|SweatGlandAdenocarcinoma|8401/3|ApocrineAdenocarcinoma
C440-C449|Skin|840|SweatGlandAdenocarcinoma|8402/3|SweatGlandAdenocarcinoma
C440-C449|Skin|840|SweatGlandAdenocarcinoma|8403/3|Spiradenocarcinoma
C440-C449|Skin|840|SweatGlandAdenocarcinoma|8407/3|MicrocysticAdnexalCarcinoma
C440-C449|Skin|840|SweatGlandAdenocarcinoma|8408/3|DigitalPapillaryEccrineCarcinoma
C440-C449|Skin|840|SweatGlandAdenocarcinoma|8409/3|EccrinePorocarcinoma
C440-C449|Skin|841|EccrineAdenocarcinoma|8410/3|SebaceousAdenocarcinoma
C440-C449|Skin|841|EccrineAdenocarcinoma|8413/3|EccrineAdenocarcinoma
C440-C449|Skin|842|CeruminousAdenocarcinoma|8420/3|CeruminousAdenocarcinoma
C440-C449|Skin|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C440-C449|Skin|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C440-C449|Skin|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C440-C449|Skin|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C440-C449|Skin|854|PagetDiseaseExtramammary|8542/3|PagetDiseaseExtramammary
C440-C449|Skin|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C440-C449|Skin|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C440-C449|Skin|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C440-C449|Skin|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C440-C449|Skin|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C440-C449|Skin|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C440-C449|Skin|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C440-C449|Skin|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C440-C449|Skin|872|Melanoma|8720/2|Stage0SkinMelanoma
C440-C449|Skin|872|Melanoma|8720/3|Melanoma
C440-C449|Skin|872|Melanoma|8721/3|NodularMelanoma
C440-C449|Skin|872|Melanoma|8722/3|BalloonCellMelanoma
C440-C449|Skin|872|Melanoma|8723/3|RegressingMelanoma
C440-C449|Skin|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C440-C449|Skin|874|Nevus|8740/3|MelanomaInJunctionalNevus
C440-C449|Skin|874|Nevus|8741/2|PrecancerousMelanosis
C440-C449|Skin|874|Nevus|8741/3|Melanoma
C440-C449|Skin|874|Nevus|8742/2|LentigoMaligna
C440-C449|Skin|874|Nevus|8742/3|LentigoMalignaMelanoma
C440-C449|Skin|874|Nevus|8743/2|SuperficialSpreadingMelanoma
C440-C449|Skin|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C440-C449|Skin|874|Nevus|8744/3|AcralLentiginousMelanoma
C440-C449|Skin|874|Nevus|8745/3|DesmoplasticMelanoma
C440-C449|Skin|874|Nevus|8746/3|MucosalLentiginousMelanoma
C440-C449|Skin|876|Nevus|8761/3|GiantCongenitalNevus
C440-C449|Skin|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C440-C449|Skin|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C440-C449|Skin|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C440-C449|Skin|878|MelanomaArisingFromBlueNevus|8780/3|MelanomaArisingFromBlueNevus
C440-C449|Skin|880|Sarcoma|8800/3|Sarcoma
C440-C449|Skin|880|Sarcoma|8801/3|SpindleCellSarcoma
C440-C449|Skin|880|Sarcoma|8802/3|GiantCellSarcoma
C440-C449|Skin|880|Sarcoma|8803/3|SmallCellSarcoma
C440-C449|Skin|880|Sarcoma|8804/3|SarcomaEpithelioid
C440-C449|Skin|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C440-C449|Skin|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C440-C449|Skin|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C440-C449|Skin|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C440-C449|Skin|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C440-C449|Skin|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C440-C449|Skin|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C440-C449|Skin|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C440-C449|Skin|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C440-C449|Skin|883|BenignFibrousHistiocytoma|8832/3|DermatofibrosarcomaProtuberans
C440-C449|Skin|883|BenignFibrousHistiocytoma|8833/3|DermatofibrosarcomaProtuberans
C440-C449|Skin|885|Liposarcoma|8850/3|Liposarcoma
C440-C449|Skin|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C440-C449|Skin|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C440-C449|Skin|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C440-C449|Skin|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C440-C449|Skin|885|Liposarcoma|8855/3|Liposarcoma
C440-C449|Skin|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C440-C449|Skin|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C440-C449|Skin|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C440-C449|Skin|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C440-C449|Skin|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C440-C449|Skin|889|MyomatousNeoplasm|8895/3|Myosarcoma
C440-C449|Skin|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C440-C449|Skin|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C440-C449|Skin|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C440-C449|Skin|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C440-C449|Skin|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C440-C449|Skin|898|Carcinosarcoma|8980/3|Carcinosarcoma
C440-C449|Skin|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C440-C449|Skin|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C440-C449|Skin|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C440-C449|Skin|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C440-C449|Skin|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C440-C449|Skin|914|KaposiSarcoma|9140/3|KaposiSarcoma
C440-C449|Skin|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C440-C449|Skin|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C440-C449|Skin|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C440-C449|Skin|959|Lymphoma|9590/3|Lymphoma
C440-C449|Skin|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C440-C449|Skin|959|Lymphoma|9596/3|CompositeLymphoma
C440-C449|Skin|959|Lymphoma|9597/3|CrostisDisease
C440-C449|Skin|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C440-C449|Skin|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C440-C449|Skin|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C440-C449|Skin|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C440-C449|Skin|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C440-C449|Skin|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C440-C449|Skin|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C440-C449|Skin|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C440-C449|Skin|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C440-C449|Skin|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C440-C449|Skin|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C440-C449|Skin|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C440-C449|Skin|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C440-C449|Skin|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C440-C449|Skin|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C440-C449|Skin|967|BCellLymphomas|9673/3|MantleCellLymphoma
C440-C449|Skin|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C440-C449|Skin|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C440-C449|Skin|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C440-C449|Skin|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C440-C449|Skin|969|FollicularAdenoma|9690/3|LymphomaFollicular
C440-C449|Skin|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C440-C449|Skin|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C440-C449|Skin|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C440-C449|Skin|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C440-C449|Skin|970|TCellLymphoma|9700/3|MycosisFungoides
C440-C449|Skin|970|TCellLymphoma|9701/3|SezarySyndrome
C440-C449|Skin|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C440-C449|Skin|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C440-C449|Skin|970|TCellLymphoma|9708/3|TCellLymphoma
C440-C449|Skin|970|TCellLymphoma|9709/3|CutaneousTCellNonHodgkinLymphoma
C440-C449|Skin|971|AdultNonHodgkinLymphoma|9718/3|CALCL
C440-C449|Skin|972|LymphoblasticLymphoma|9725/3|HydroaVacciniformeLikeLymphoma
C440-C449|Skin|972|LymphoblasticLymphoma|9726/3|TCellLymphoma
C440-C449|Skin|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C440-C449|Skin|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C440-C449|Skin|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C440-C449|Skin|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C440-C449|Skin|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C440-C449|Skin|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C470-C476,C478-C479|PeripheralNerve|868|Paraganglioma|8680/3|MalignantParaganglioma
C470-C476,C478-C479|PeripheralNerve|869|MalignantExtraAdrenalParaganglioma|8693/3|MalignantExtraAdrenalParaganglioma
C470-C476,C478-C479|PeripheralNerve|880|Sarcoma|8800/3|Sarcoma
C470-C476,C478-C479|PeripheralNerve|880|Sarcoma|8801/3|SpindleCellSarcoma
C470-C476,C478-C479|PeripheralNerve|880|Sarcoma|8802/3|GiantCellSarcoma
C470-C476,C478-C479|PeripheralNerve|880|Sarcoma|8803/3|SmallCellSarcoma
C470-C476,C478-C479|PeripheralNerve|880|Sarcoma|8804/3|SarcomaEpithelioid
C470-C476,C478-C479|PeripheralNerve|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C470-C476,C478-C479|PeripheralNerve|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C470-C476,C478-C479|PeripheralNerve|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C470-C476,C478-C479|PeripheralNerve|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C470-C476,C478-C479|PeripheralNerve|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C470-C476,C478-C479|PeripheralNerve|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C470-C476,C478-C479|PeripheralNerve|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C470-C476,C478-C479|PeripheralNerve|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C470-C476,C478-C479|PeripheralNerve|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C470-C476,C478-C479|PeripheralNerve|883|BenignFibrousHistiocytoma|8832/3|DermatofibrosarcomaProtuberans
C470-C476,C478-C479|PeripheralNerve|883|BenignFibrousHistiocytoma|8833/3|DermatofibrosarcomaProtuberans
C470-C476,C478-C479|PeripheralNerve|884|Myxosarcoma|8840/3|Myxosarcoma
C470-C476,C478-C479|PeripheralNerve|885|Liposarcoma|8850/3|Liposarcoma
C470-C476,C478-C479|PeripheralNerve|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C470-C476,C478-C479|PeripheralNerve|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C470-C476,C478-C479|PeripheralNerve|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C470-C476,C478-C479|PeripheralNerve|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C470-C476,C478-C479|PeripheralNerve|885|Liposarcoma|8855/3|Liposarcoma
C470-C476,C478-C479|PeripheralNerve|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C470-C476,C478-C479|PeripheralNerve|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C470-C476,C478-C479|PeripheralNerve|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C470-C476,C478-C479|PeripheralNerve|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C470-C476,C478-C479|PeripheralNerve|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C470-C476,C478-C479|PeripheralNerve|889|MyomatousNeoplasm|8895/3|Myosarcoma
C470-C476,C478-C479|PeripheralNerve|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C470-C476,C478-C479|PeripheralNerve|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C470-C476,C478-C479|PeripheralNerve|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C470-C476,C478-C479|PeripheralNerve|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C470-C476,C478-C479|PeripheralNerve|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C470-C476,C478-C479|PeripheralNerve|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C470-C476,C478-C479|PeripheralNerve|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C470-C476,C478-C479|PeripheralNerve|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C470-C476,C478-C479|PeripheralNerve|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C470-C476,C478-C479|PeripheralNerve|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C470-C476,C478-C479|PeripheralNerve|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C470-C476,C478-C479|PeripheralNerve|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C470-C476,C478-C479|PeripheralNerve|904|SynovialSarcoma|9040/3|SynovialSarcoma
C470-C476,C478-C479|PeripheralNerve|904|SynovialSarcoma|9041/3|SpindleCellSynovialSarcoma
C470-C476,C478-C479|PeripheralNerve|904|SynovialSarcoma|9042/3|EpithelialSynovialSarcoma
C470-C476,C478-C479|PeripheralNerve|904|SynovialSarcoma|9043/3|BiphasicSynovialSarcoma
C470-C476,C478-C479|PeripheralNerve|904|SynovialSarcoma|9044/3|ClearCellSarcomaOfSoftTissueC0206651
C470-C476,C478-C479|PeripheralNerve|908|Teratoma|9080/3|ImmatureTeratoma
C470-C476,C478-C479|PeripheralNerve|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C470-C476,C478-C479|PeripheralNerve|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C470-C476,C478-C479|PeripheralNerve|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C470-C476,C478-C479|PeripheralNerve|908|Teratoma|9084/3|Teratoma
C470-C476,C478-C479|PeripheralNerve|908|Teratoma|9085/3|MixedGermCellTumor
C470-C476,C478-C479|PeripheralNerve|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C470-C476,C478-C479|PeripheralNerve|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C470-C476,C478-C479|PeripheralNerve|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C470-C476,C478-C479|PeripheralNerve|914|KaposiSarcoma|9140/3|KaposiSarcoma
C470-C476,C478-C479|PeripheralNerve|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C470-C476,C478-C479|PeripheralNerve|917|Lymphangiosarcoma|9170/3|Lymphangiosarcoma
C470-C476,C478-C479|PeripheralNerve|924|OsseousAndChondromatousNeoplasms|9240/3|MesenchymalChondrosarcoma
C470-C476,C478-C479|PeripheralNerve|924|OsseousAndChondromatousNeoplasms|9242/3|ClearCellChondrosarcoma
C470-C476,C478-C479|PeripheralNerve|924|OsseousAndChondromatousNeoplasms|9243/3|DedifferentiatedChondrosarcoma
C470-C476,C478-C479|PeripheralNerve|925|BoneNeoplasm|9251/3|GiantCellTumorOfSoftTissue
C470-C476,C478-C479|PeripheralNerve|925|BoneNeoplasm|9252/3|MalignantTenosynovialGiantCellTumor
C470-C476,C478-C479|PeripheralNerve|936|NeuroepitheliomaPeripheral|9364/3|NeuroepitheliomaPeripheral
C470-C476,C478-C479|PeripheralNerve|936|NeuroepitheliomaPeripheral|9365/3|AskinTumor
C470-C476,C478-C479|PeripheralNerve|937|Chordoma|9370/3|Chordoma
C470-C476,C478-C479|PeripheralNerve|937|Chordoma|9371/3|ChondroidChordoma
C470-C476,C478-C479|PeripheralNerve|937|Chordoma|9372/3|DedifferentiatedChordoma
C470-C476,C478-C479|PeripheralNerve|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C470-C476,C478-C479|PeripheralNerve|950|Neuroblastoma|9500/3|Neuroblastoma
C470-C476,C478-C479|PeripheralNerve|950|Neuroblastoma|9501/3|Medulloepithelioma
C470-C476,C478-C479|PeripheralNerve|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C470-C476,C478-C479|PeripheralNerve|950|Neuroblastoma|9503/3|Neuroepithelioma
C470-C476,C478-C479|PeripheralNerve|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C470-C476,C478-C479|PeripheralNerve|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C470-C476,C478-C479|PeripheralNerve|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C470-C476,C478-C479|PeripheralNerve|954|MalignantPeripheralNerveSheathTumor|9542/3|MalignantPeripheralNerveSheathTumor
C470-C476,C478-C479|PeripheralNerve|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C470-C476,C478-C479|PeripheralNerve|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C470-C476,C478-C479|PeripheralNerve|957|Perineurioma|9571/3|MalignantPerineurioma
C470-C476,C478-C479|PeripheralNerve|958|GranularCellTumor|9580/3|MalignantGranularCellTumor
C470-C476,C478-C479|PeripheralNerve|958|GranularCellTumor|9581/3|AlveolarSoftPartSarcoma
C470-C476,C478-C479|PeripheralNerve|959|Lymphoma|9590/3|Lymphoma
C470-C476,C478-C479|PeripheralNerve|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C470-C476,C478-C479|PeripheralNerve|959|Lymphoma|9596/3|CompositeLymphoma
C470-C476,C478-C479|PeripheralNerve|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C470-C476,C478-C479|PeripheralNerve|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C470-C476,C478-C479|PeripheralNerve|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C470-C476,C478-C479|PeripheralNerve|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C470-C476,C478-C479|PeripheralNerve|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C470-C476,C478-C479|PeripheralNerve|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C470-C476,C478-C479|PeripheralNerve|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C470-C476,C478-C479|PeripheralNerve|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C470-C476,C478-C479|PeripheralNerve|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C470-C476,C478-C479|PeripheralNerve|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C470-C476,C478-C479|PeripheralNerve|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C470-C476,C478-C479|PeripheralNerve|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C470-C476,C478-C479|PeripheralNerve|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C470-C476,C478-C479|PeripheralNerve|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C470-C476,C478-C479|PeripheralNerve|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C470-C476,C478-C479|PeripheralNerve|967|BCellLymphomas|9673/3|MantleCellLymphoma
C470-C476,C478-C479|PeripheralNerve|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C470-C476,C478-C479|PeripheralNerve|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C470-C476,C478-C479|PeripheralNerve|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C470-C476,C478-C479|PeripheralNerve|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C470-C476,C478-C479|PeripheralNerve|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C470-C476,C478-C479|PeripheralNerve|969|FollicularAdenoma|9690/3|LymphomaFollicular
C470-C476,C478-C479|PeripheralNerve|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C470-C476,C478-C479|PeripheralNerve|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C470-C476,C478-C479|PeripheralNerve|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C470-C476,C478-C479|PeripheralNerve|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C470-C476,C478-C479|PeripheralNerve|970|TCellLymphoma|9701/3|SezarySyndrome
C470-C476,C478-C479|PeripheralNerve|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C470-C476,C478-C479|PeripheralNerve|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C470-C476,C478-C479|PeripheralNerve|970|TCellLymphoma|9708/3|TCellLymphoma
C470-C476,C478-C479|PeripheralNerve|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C470-C476,C478-C479|PeripheralNerve|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C470-C476,C478-C479|PeripheralNerve|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C470-C476,C478-C479|PeripheralNerve|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C470-C476,C478-C479|PeripheralNerve|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C470-C476,C478-C479|PeripheralNerve|972|LymphoblasticLymphoma|9726/3|TCellLymphoma
C470-C476,C478-C479|PeripheralNerve|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C470-C476,C478-C479|PeripheralNerve|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C470-C476,C478-C479|PeripheralNerve|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C470-C476,C478-C479|PeripheralNerve|973|Plasmacytoma|9731/3|Plasmacytoma
C470-C476,C478-C479|PeripheralNerve|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C470-C476,C478-C479|PeripheralNerve|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C470-C476,C478-C479|PeripheralNerve|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C470-C476,C478-C479|PeripheralNerve|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C470-C476,C478-C479|PeripheralNerve|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C470-C476,C478-C479|PeripheralNerve|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C470-C476,C478-C479|PeripheralNerve|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C470-C476,C478-C479|PeripheralNerve|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C470-C476,C478-C479|PeripheralNerve|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C470-C476,C478-C479|PeripheralNerve|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C470-C476,C478-C479|PeripheralNerve|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C470-C476,C478-C479|PeripheralNerve|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C470-C476,C478-C479|PeripheralNerve|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C470-C476,C478-C479|PeripheralNerve|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C470-C476,C478-C479|PeripheralNerve|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C470-C476,C478-C479|PeripheralNerve|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9812/3|null
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9813/3|null
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9814/3|null
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9817/3|null
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9818/3|null
C470-C476,C478-C479|PeripheralNerve|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C470-C476,C478-C479|PeripheralNerve|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C470-C476,C478-C479|PeripheralNerve|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C470-C476,C478-C479|PeripheralNerve|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C470-C476,C478-C479|PeripheralNerve|993|MyeloidSarcoma|9930/3|MyeloidSarcoma
C470-C476,C478-C479|PeripheralNerve|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C470-C476,C478-C479|PeripheralNerve|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C470-C476,C478-C479|PeripheralNerve|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C470-C476,C478-C479|PeripheralNerve|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C480-C482,C488|RetroperitonealSpace|846|PapillarySerousCystadenocarcinoma|8461/3|SerousSurfacePapillaryCarcinoma
C480-C482,C488|RetroperitonealSpace|868|Paraganglioma|8680/3|MalignantParaganglioma
C480-C482,C488|RetroperitonealSpace|869|MalignantExtraAdrenalParaganglioma|8693/3|MalignantExtraAdrenalParaganglioma
C480-C482,C488|RetroperitonealSpace|871|MalignantGlomusTumor|8714/3|MalignantPEComa
C480-C482,C488|RetroperitonealSpace|880|Sarcoma|8800/3|Sarcoma
C480-C482,C488|RetroperitonealSpace|880|Sarcoma|8801/3|SpindleCellSarcoma
C480-C482,C488|RetroperitonealSpace|880|Sarcoma|8802/3|GiantCellSarcoma
C480-C482,C488|RetroperitonealSpace|880|Sarcoma|8803/3|SmallCellSarcoma
C480-C482,C488|RetroperitonealSpace|880|Sarcoma|8804/3|SarcomaEpithelioid
C480-C482,C488|RetroperitonealSpace|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C480-C482,C488|RetroperitonealSpace|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C480-C482,C488|RetroperitonealSpace|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C480-C482,C488|RetroperitonealSpace|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C480-C482,C488|RetroperitonealSpace|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C480-C482,C488|RetroperitonealSpace|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C480-C482,C488|RetroperitonealSpace|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C480-C482,C488|RetroperitonealSpace|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C480-C482,C488|RetroperitonealSpace|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C480-C482,C488|RetroperitonealSpace|884|Myxosarcoma|8840/3|Myxosarcoma
C480-C482,C488|RetroperitonealSpace|885|Liposarcoma|8850/3|Liposarcoma
C480-C482,C488|RetroperitonealSpace|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C480-C482,C488|RetroperitonealSpace|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C480-C482,C488|RetroperitonealSpace|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C480-C482,C488|RetroperitonealSpace|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C480-C482,C488|RetroperitonealSpace|885|Liposarcoma|8855/3|Liposarcoma
C480-C482,C488|RetroperitonealSpace|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C480-C482,C488|RetroperitonealSpace|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C480-C482,C488|RetroperitonealSpace|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C480-C482,C488|RetroperitonealSpace|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C480-C482,C488|RetroperitonealSpace|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C480-C482,C488|RetroperitonealSpace|889|MyomatousNeoplasm|8895/3|Myosarcoma
C480-C482,C488|RetroperitonealSpace|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C480-C482,C488|RetroperitonealSpace|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C480-C482,C488|RetroperitonealSpace|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C480-C482,C488|RetroperitonealSpace|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C480-C482,C488|RetroperitonealSpace|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C480-C482,C488|RetroperitonealSpace|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C480-C482,C488|RetroperitonealSpace|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C480-C482,C488|RetroperitonealSpace|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C480-C482,C488|RetroperitonealSpace|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C480-C482,C488|RetroperitonealSpace|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C480-C482,C488|RetroperitonealSpace|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C480-C482,C488|RetroperitonealSpace|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C480-C482,C488|RetroperitonealSpace|905|MalignantMesothelioma|9050/3|MalignantMesothelioma
C480-C482,C488|RetroperitonealSpace|905|MalignantMesothelioma|9051/3|SarcomatoidMesothelioma
C480-C482,C488|RetroperitonealSpace|905|MalignantMesothelioma|9052/3|Mesothelioma
C480-C482,C488|RetroperitonealSpace|905|MalignantMesothelioma|9053/3|BiphasicMesothelioma
C480-C482,C488|RetroperitonealSpace|906|GermCellTumor|9060/3|Dysgerminoma
C480-C482,C488|RetroperitonealSpace|906|GermCellTumor|9064/3|Germinoma
C480-C482,C488|RetroperitonealSpace|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C480-C482,C488|RetroperitonealSpace|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C480-C482,C488|RetroperitonealSpace|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C480-C482,C488|RetroperitonealSpace|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C480-C482,C488|RetroperitonealSpace|908|Teratoma|9080/3|ImmatureTeratoma
C480-C482,C488|RetroperitonealSpace|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C480-C482,C488|RetroperitonealSpace|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C480-C482,C488|RetroperitonealSpace|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C480-C482,C488|RetroperitonealSpace|908|Teratoma|9084/3|Teratoma
C480-C482,C488|RetroperitonealSpace|908|Teratoma|9085/3|MixedGermCellTumor
C480-C482,C488|RetroperitonealSpace|911|Mesonephroma|9110/3|Mesonephroma
C480-C482,C488|RetroperitonealSpace|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C480-C482,C488|RetroperitonealSpace|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C480-C482,C488|RetroperitonealSpace|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C480-C482,C488|RetroperitonealSpace|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C480-C482,C488|RetroperitonealSpace|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C480-C482,C488|RetroperitonealSpace|950|Neuroblastoma|9500/3|Neuroblastoma
C480-C482,C488|RetroperitonealSpace|950|Neuroblastoma|9501/3|Medulloepithelioma
C480-C482,C488|RetroperitonealSpace|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C480-C482,C488|RetroperitonealSpace|950|Neuroblastoma|9503/3|Neuroepithelioma
C480-C482,C488|RetroperitonealSpace|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C480-C482,C488|RetroperitonealSpace|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C480-C482,C488|RetroperitonealSpace|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C480-C482,C488|RetroperitonealSpace|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C480-C482,C488|RetroperitonealSpace|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C480-C482,C488|RetroperitonealSpace|957|Perineurioma|9571/3|MalignantPerineurioma
C480-C482,C488|RetroperitonealSpace|959|Lymphoma|9590/3|Lymphoma
C480-C482,C488|RetroperitonealSpace|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C480-C482,C488|RetroperitonealSpace|959|Lymphoma|9596/3|CompositeLymphoma
C480-C482,C488|RetroperitonealSpace|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C480-C482,C488|RetroperitonealSpace|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C480-C482,C488|RetroperitonealSpace|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C480-C482,C488|RetroperitonealSpace|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C480-C482,C488|RetroperitonealSpace|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C480-C482,C488|RetroperitonealSpace|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C480-C482,C488|RetroperitonealSpace|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C480-C482,C488|RetroperitonealSpace|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C480-C482,C488|RetroperitonealSpace|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C480-C482,C488|RetroperitonealSpace|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C480-C482,C488|RetroperitonealSpace|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C480-C482,C488|RetroperitonealSpace|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C480-C482,C488|RetroperitonealSpace|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C480-C482,C488|RetroperitonealSpace|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C480-C482,C488|RetroperitonealSpace|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C480-C482,C488|RetroperitonealSpace|967|BCellLymphomas|9673/3|MantleCellLymphoma
C480-C482,C488|RetroperitonealSpace|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C480-C482,C488|RetroperitonealSpace|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C480-C482,C488|RetroperitonealSpace|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C480-C482,C488|RetroperitonealSpace|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C480-C482,C488|RetroperitonealSpace|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C480-C482,C488|RetroperitonealSpace|969|FollicularAdenoma|9690/3|LymphomaFollicular
C480-C482,C488|RetroperitonealSpace|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C480-C482,C488|RetroperitonealSpace|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C480-C482,C488|RetroperitonealSpace|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C480-C482,C488|RetroperitonealSpace|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C480-C482,C488|RetroperitonealSpace|970|TCellLymphoma|9701/3|SezarySyndrome
C480-C482,C488|RetroperitonealSpace|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C480-C482,C488|RetroperitonealSpace|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C480-C482,C488|RetroperitonealSpace|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C480-C482,C488|RetroperitonealSpace|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C480-C482,C488|RetroperitonealSpace|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C480-C482,C488|RetroperitonealSpace|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C480-C482,C488|RetroperitonealSpace|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C480-C482,C488|RetroperitonealSpace|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C480-C482,C488|RetroperitonealSpace|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C480-C482,C488|RetroperitonealSpace|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C480-C482,C488|RetroperitonealSpace|973|Plasmacytoma|9731/3|Plasmacytoma
C480-C482,C488|RetroperitonealSpace|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C480-C482,C488|RetroperitonealSpace|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C480-C482,C488|RetroperitonealSpace|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C480-C482,C488|RetroperitonealSpace|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C480-C482,C488|RetroperitonealSpace|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C480-C482,C488|RetroperitonealSpace|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C480-C482,C488|RetroperitonealSpace|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C480-C482,C488|RetroperitonealSpace|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C480-C482,C488|RetroperitonealSpace|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C480-C482,C488|RetroperitonealSpace|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C480-C482,C488|RetroperitonealSpace|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C480-C482,C488|RetroperitonealSpace|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C480-C482,C488|RetroperitonealSpace|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C480-C482,C488|RetroperitonealSpace|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C480-C482,C488|RetroperitonealSpace|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C480-C482,C488|RetroperitonealSpace|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9812/3|null
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9813/3|null
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9814/3|null
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9817/3|null
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9818/3|null
C480-C482,C488|RetroperitonealSpace|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C480-C482,C488|RetroperitonealSpace|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C480-C482,C488|RetroperitonealSpace|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C480-C482,C488|RetroperitonealSpace|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C480-C482,C488|RetroperitonealSpace|993|MyeloidSarcoma|9930/3|MyeloidSarcoma
C480-C482,C488|RetroperitonealSpace|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C480-C482,C488|RetroperitonealSpace|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C480-C482,C488|RetroperitonealSpace|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C480-C482,C488|RetroperitonealSpace|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C500-C506,C508-C509|Breast|801|Carcinoma|8010/2|InSituCancer
C500-C506,C508-C509|Breast|801|Carcinoma|8010/3|CarcinomaNOSDNE
C500-C506,C508-C509|Breast|801|Carcinoma|8011/3|MalignantEpithelioma
C500-C506,C508-C509|Breast|801|Carcinoma|8012/3|LargeCellCarcinoma
C500-C506,C508-C509|Breast|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C500-C506,C508-C509|Breast|801|Carcinoma|8014/3|LargeCellCarcinoma
C500-C506,C508-C509|Breast|801|Carcinoma|8015/3|GlassyCellCarcinoma
C500-C506,C508-C509|Breast|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C500-C506,C508-C509|Breast|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C500-C506,C508-C509|Breast|802|Carcinoma|8022/3|PleomorphicCarcinoma
C500-C506,C508-C509|Breast|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C500-C506,C508-C509|Breast|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C500-C506,C508-C509|Breast|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C500-C506,C508-C509|Breast|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C500-C506,C508-C509|Breast|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C500-C506,C508-C509|Breast|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C500-C506,C508-C509|Breast|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C500-C506,C508-C509|Breast|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C500-C506,C508-C509|Breast|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C500-C506,C508-C509|Breast|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C500-C506,C508-C509|Breast|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C500-C506,C508-C509|Breast|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C500-C506,C508-C509|Breast|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C500-C506,C508-C509|Breast|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C500-C506,C508-C509|Breast|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8140/3|Adenocarcinoma
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C500-C506,C508-C509|Breast|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C500-C506,C508-C509|Breast|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C500-C506,C508-C509|Breast|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C500-C506,C508-C509|Breast|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C500-C506,C508-C509|Breast|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C500-C506,C508-C509|Breast|823|SolidCarcinoma|8230/2|InSituCancer
C500-C506,C508-C509|Breast|823|SolidCarcinoma|8230/3|SolidCarcinoma
C500-C506,C508-C509|Breast|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C500-C506,C508-C509|Breast|825|BronchioloalveolarAdenocarcinoma|8251/3|BronchioloalveolarAdenocarcinoma
C500-C506,C508-C509|Breast|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C500-C506,C508-C509|Breast|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C500-C506,C508-C509|Breast|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C500-C506,C508-C509|Breast|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C500-C506,C508-C509|Breast|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C500-C506,C508-C509|Breast|831|ClearCellAdenocarcinoma|8314/3|LipidRichCarcinoma
C500-C506,C508-C509|Breast|831|ClearCellAdenocarcinoma|8315/3|GlycogenRichCarcinoma
C500-C506,C508-C509|Breast|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C500-C506,C508-C509|Breast|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C500-C506,C508-C509|Breast|840|SweatGlandAdenocarcinoma|8401/3|ApocrineAdenocarcinoma
C500-C506,C508-C509|Breast|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C500-C506,C508-C509|Breast|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C500-C506,C508-C509|Breast|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C500-C506,C508-C509|Breast|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8500/1|DuctalCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8500/2|DuctalBreastCarcinomaInSitu
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8500/3|InvasiveBreastCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8501/2|Comedocarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8501/3|Comedocarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8502/3|SecretoryBreastCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8503/2|IntraductalPapillaryBreastCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8503/3|IntraductalPapillaryBreastCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8504/2|IntracysticPapillaryBreastCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8504/3|IntracysticPapillaryBreastCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8507/2|MicropapillaryCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8507/3|MicropapillaryCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8508/3|SecretoryBreastCarcinoma
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8509/2|SolidPapillaryCarcinomaInSitu
C500-C506,C508-C509|Breast|850|DuctalCarcinoma|8509/3|PapillaryCarcinoma
C500-C506,C508-C509|Breast|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C500-C506,C508-C509|Breast|851|MedullaryCarcinoma|8512/3|MedullaryCarcinoma
C500-C506,C508-C509|Breast|851|MedullaryCarcinoma|8513/3|MedullaryCarcinoma
C500-C506,C508-C509|Breast|851|MedullaryCarcinoma|8514/3|DesmoplasticNodularMedulloblastoma
C500-C506,C508-C509|Breast|851|MedullaryCarcinoma|8519/2|PleomorphicLobularCarcinomaInSitu
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8520/2|LobularBreastCarcinomaInSitu
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8520/3|CarcinomaLobular
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8521/3|InvasiveDuctalBreastCarcinoma
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8522/2|BreastCarcinoma
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8522/3|IntraductalAndLobularCarcinoma
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8523/2|InfiltratingDuctAndTubularCarcinoma
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8523/3|InfiltratingDuctAndTubularCarcinoma
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8524/3|InvasiveLobularBreastCarcinoma
C500-C506,C508-C509|Breast|852|IntraductalAndLobularCarcinoma|8525/3|TerminalDuctAdenocarcinoma
C500-C506,C508-C509|Breast|853|InflammatoryCarcinoma|8530/3|InflammatoryCarcinoma
C500-C506,C508-C509|Breast|854|PagetsDiseaseMammary|8540/3|PagetsDiseaseMammary
C500-C506,C508-C509|Breast|854|PagetsDiseaseMammary|8541/3|PagetsDiseaseMammary
C500-C506,C508-C509|Breast|854|PagetsDiseaseMammary|8543/3|PagetDisease
C500-C506,C508-C509|Breast|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C500-C506,C508-C509|Breast|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C500-C506,C508-C509|Breast|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C500-C506,C508-C509|Breast|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C500-C506,C508-C509|Breast|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C500-C506,C508-C509|Breast|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C500-C506,C508-C509|Breast|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C500-C506,C508-C509|Breast|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C500-C506,C508-C509|Breast|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C500-C506,C508-C509|Breast|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C500-C506,C508-C509|Breast|880|Sarcoma|8800/3|Sarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8801/3|SpindleCellSarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8802/3|GiantCellSarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8803/3|SmallCellSarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8804/3|SarcomaEpithelioid
C500-C506,C508-C509|Breast|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C500-C506,C508-C509|Breast|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C500-C506,C508-C509|Breast|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C500-C506,C508-C509|Breast|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C500-C506,C508-C509|Breast|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C500-C506,C508-C509|Breast|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C500-C506,C508-C509|Breast|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8850/3|Liposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C500-C506,C508-C509|Breast|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8855/3|Liposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C500-C506,C508-C509|Breast|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C500-C506,C508-C509|Breast|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C500-C506,C508-C509|Breast|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C500-C506,C508-C509|Breast|889|MyomatousNeoplasm|8895/3|Myosarcoma
C500-C506,C508-C509|Breast|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C500-C506,C508-C509|Breast|893|StromalSarcoma|8935/3|StromalSarcoma
C500-C506,C508-C509|Breast|898|Carcinosarcoma|8980/3|Carcinosarcoma
C500-C506,C508-C509|Breast|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C500-C506,C508-C509|Breast|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C500-C506,C508-C509|Breast|898|Carcinosarcoma|8983/3|AdenomyoepitheliomaWithCarcinoma
C500-C506,C508-C509|Breast|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C500-C506,C508-C509|Breast|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C500-C506,C508-C509|Breast|902|PhyllodesTumor|9020/3|MalignantPhyllodesTumor
C500-C506,C508-C509|Breast|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C500-C506,C508-C509|Breast|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C500-C506,C508-C509|Breast|913|Hemangioendothelioma|9133/3|EpithelioidHemangioendothelioma
C500-C506,C508-C509|Breast|958|GranularCellTumor|9580/3|MalignantGranularCellTumor
C500-C506,C508-C509|Breast|958|GranularCellTumor|9581/3|AlveolarSoftPartSarcoma
C500-C506,C508-C509|Breast|959|Lymphoma|9590/3|Lymphoma
C500-C506,C508-C509|Breast|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C500-C506,C508-C509|Breast|959|Lymphoma|9596/3|CompositeLymphoma
C500-C506,C508-C509|Breast|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C500-C506,C508-C509|Breast|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C500-C506,C508-C509|Breast|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C500-C506,C508-C509|Breast|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C500-C506,C508-C509|Breast|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C500-C506,C508-C509|Breast|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C500-C506,C508-C509|Breast|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C500-C506,C508-C509|Breast|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C500-C506,C508-C509|Breast|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C500-C506,C508-C509|Breast|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C500-C506,C508-C509|Breast|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C500-C506,C508-C509|Breast|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C500-C506,C508-C509|Breast|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C500-C506,C508-C509|Breast|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C500-C506,C508-C509|Breast|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C500-C506,C508-C509|Breast|967|BCellLymphomas|9673/3|MantleCellLymphoma
C500-C506,C508-C509|Breast|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C500-C506,C508-C509|Breast|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C500-C506,C508-C509|Breast|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C500-C506,C508-C509|Breast|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C500-C506,C508-C509|Breast|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C500-C506,C508-C509|Breast|969|FollicularAdenoma|9690/3|LymphomaFollicular
C500-C506,C508-C509|Breast|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C500-C506,C508-C509|Breast|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C500-C506,C508-C509|Breast|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C500-C506,C508-C509|Breast|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C500-C506,C508-C509|Breast|970|TCellLymphoma|9701/3|SezarySyndrome
C500-C506,C508-C509|Breast|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C500-C506,C508-C509|Breast|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C500-C506,C508-C509|Breast|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C500-C506,C508-C509|Breast|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C500-C506,C508-C509|Breast|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C500-C506,C508-C509|Breast|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C500-C506,C508-C509|Breast|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C500-C506,C508-C509|Breast|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C500-C506,C508-C509|Breast|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C500-C506,C508-C509|Breast|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C500-C506,C508-C509|Breast|973|Plasmacytoma|9731/3|Plasmacytoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C500-C506,C508-C509|Breast|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C500-C506,C508-C509|Breast|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C500-C506,C508-C509|Breast|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C500-C506,C508-C509|Breast|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C500-C506,C508-C509|Breast|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C500-C506,C508-C509|Breast|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C500-C506,C508-C509|Breast|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C500-C506,C508-C509|Breast|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C500-C506,C508-C509|Breast|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C500-C506,C508-C509|Breast|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C500-C506,C508-C509|Breast|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C500-C506,C508-C509|Breast|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9812/3|null
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9813/3|null
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9814/3|null
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9817/3|null
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9818/3|null
C500-C506,C508-C509|Breast|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C500-C506,C508-C509|Breast|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C500-C506,C508-C509|Breast|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C500-C506,C508-C509|Breast|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C500-C506,C508-C509|Breast|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C500-C506,C508-C509|Breast|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C500-C506,C508-C509|Breast|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C500-C506,C508-C509|Breast|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C510-C512,C518, C529|Vagina|801|Carcinoma|8010/2|InSituCancer
C510-C512,C518, C529|Vagina|801|Carcinoma|8010/3|CarcinomaNOSDNE
C510-C512,C518, C529|Vagina|801|Carcinoma|8011/3|MalignantEpithelioma
C510-C512,C518, C529|Vagina|801|Carcinoma|8012/3|LargeCellCarcinoma
C510-C512,C518, C529|Vagina|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C510-C512,C518, C529|Vagina|801|Carcinoma|8014/3|LargeCellCarcinoma
C510-C512,C518, C529|Vagina|801|Carcinoma|8015/3|GlassyCellCarcinoma
C510-C512,C518, C529|Vagina|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C510-C512,C518, C529|Vagina|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C510-C512,C518, C529|Vagina|802|Carcinoma|8022/3|PleomorphicCarcinoma
C510-C512,C518, C529|Vagina|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C510-C512,C518, C529|Vagina|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C510-C512,C518, C529|Vagina|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C510-C512,C518, C529|Vagina|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C510-C512,C518, C529|Vagina|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8071/2|KeratinizingSquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8077/2|IntraepithelialNeoplasia
C510-C512,C518, C529|Vagina|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C510-C512,C518, C529|Vagina|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C510-C512,C518, C529|Vagina|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C510-C512,C518, C529|Vagina|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C510-C512,C518, C529|Vagina|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C510-C512,C518, C529|Vagina|809|BasalCellCarcinoma|8090/3|BasalCellCarcinoma
C510-C512,C518, C529|Vagina|809|BasalCellCarcinoma|8091/3|SuperficialBasalCellCarcinoma
C510-C512,C518, C529|Vagina|809|BasalCellCarcinoma|8092/3|SkinInfiltratingBasalCellCarcinoma
C510-C512,C518, C529|Vagina|809|BasalCellCarcinoma|8093/3|FibroepitheliomaOfPinkus
C510-C512,C518, C529|Vagina|809|BasalCellCarcinoma|8094/3|SkinBasosquamousCellCarcinoma
C510-C512,C518, C529|Vagina|809|BasalCellCarcinoma|8095/3|SkinMetatypicalCarcinoma
C510-C512,C518, C529|Vagina|809|BasalCellCarcinoma|8097/3|SkinNodularBasalCellCarcinoma
C510-C512,C518, C529|Vagina|809|BasalCellCarcinoma|8098/3|SkinAdenoidBasalCellCarcinoma
C510-C512,C518, C529|Vagina|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C510-C512,C518, C529|Vagina|811|PilomatricalCarcinoma|8110/3|PilomatricalCarcinoma
C510-C512,C518, C529|Vagina|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C510-C512,C518, C529|Vagina|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C510-C512,C518, C529|Vagina|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C510-C512,C518, C529|Vagina|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C510-C512,C518, C529|Vagina|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C510-C512,C518, C529|Vagina|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C510-C512,C518, C529|Vagina|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C510-C512,C518, C529|Vagina|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C510-C512,C518, C529|Vagina|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8140/3|Adenocarcinoma
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C510-C512,C518, C529|Vagina|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C510-C512,C518, C529|Vagina|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C510-C512,C518, C529|Vagina|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C510-C512,C518, C529|Vagina|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C510-C512,C518, C529|Vagina|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C510-C512,C518, C529|Vagina|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C510-C512,C518, C529|Vagina|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C510-C512,C518, C529|Vagina|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C510-C512,C518, C529|Vagina|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C510-C512,C518, C529|Vagina|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C510-C512,C518, C529|Vagina|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C510-C512,C518, C529|Vagina|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C510-C512,C518, C529|Vagina|838|CarcinomaEndometrioid|8380/3|CarcinomaEndometrioid
C510-C512,C518, C529|Vagina|840|SweatGlandAdenocarcinoma|8401/3|ApocrineAdenocarcinoma
C510-C512,C518, C529|Vagina|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C510-C512,C518, C529|Vagina|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C510-C512,C518, C529|Vagina|848|MucinousAdenocarcinoma|8482/3|AdenocarcinomaEndocervicalType
C510-C512,C518, C529|Vagina|854|PagetDiseaseExtramammary|8542/3|PagetDiseaseExtramammary
C510-C512,C518, C529|Vagina|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C510-C512,C518, C529|Vagina|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C510-C512,C518, C529|Vagina|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C510-C512,C518, C529|Vagina|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C510-C512,C518, C529|Vagina|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C510-C512,C518, C529|Vagina|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C510-C512,C518, C529|Vagina|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C510-C512,C518, C529|Vagina|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C510-C512,C518, C529|Vagina|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C510-C512,C518, C529|Vagina|872|Melanoma|8720/2|Stage0SkinMelanoma
C510-C512,C518, C529|Vagina|872|Melanoma|8720/3|Melanoma
C510-C512,C518, C529|Vagina|872|Melanoma|8721/3|NodularMelanoma
C510-C512,C518, C529|Vagina|872|Melanoma|8722/3|BalloonCellMelanoma
C510-C512,C518, C529|Vagina|872|Melanoma|8723/3|RegressingMelanoma
C510-C512,C518, C529|Vagina|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C510-C512,C518, C529|Vagina|874|Nevus|8740/3|MelanomaInJunctionalNevus
C510-C512,C518, C529|Vagina|874|Nevus|8741/2|PrecancerousMelanosis
C510-C512,C518, C529|Vagina|874|Nevus|8741/3|Melanoma
C510-C512,C518, C529|Vagina|874|Nevus|8742/2|LentigoMaligna
C510-C512,C518, C529|Vagina|874|Nevus|8742/3|LentigoMalignaMelanoma
C510-C512,C518, C529|Vagina|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C510-C512,C518, C529|Vagina|874|Nevus|8745/3|DesmoplasticMelanoma
C510-C512,C518, C529|Vagina|874|Nevus|8746/3|MucosalLentiginousMelanoma
C510-C512,C518, C529|Vagina|876|Nevus|8761/3|GiantCongenitalNevus
C510-C512,C518, C529|Vagina|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C510-C512,C518, C529|Vagina|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C510-C512,C518, C529|Vagina|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8800/3|Sarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8801/3|SpindleCellSarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8802/3|GiantCellSarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8803/3|SmallCellSarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8804/3|SarcomaEpithelioid
C510-C512,C518, C529|Vagina|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C510-C512,C518, C529|Vagina|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C510-C512,C518, C529|Vagina|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C510-C512,C518, C529|Vagina|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C510-C512,C518, C529|Vagina|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C510-C512,C518, C529|Vagina|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C510-C512,C518, C529|Vagina|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C510-C512,C518, C529|Vagina|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C510-C512,C518, C529|Vagina|883|BenignFibrousHistiocytoma|8832/3|DermatofibrosarcomaProtuberans
C510-C512,C518, C529|Vagina|885|Liposarcoma|8850/3|Liposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C510-C512,C518, C529|Vagina|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8855/3|Liposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C510-C512,C518, C529|Vagina|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C510-C512,C518, C529|Vagina|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C510-C512,C518, C529|Vagina|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C510-C512,C518, C529|Vagina|889|MyomatousNeoplasm|8895/3|Myosarcoma
C510-C512,C518, C529|Vagina|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C510-C512,C518, C529|Vagina|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C510-C512,C518, C529|Vagina|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C510-C512,C518, C529|Vagina|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C510-C512,C518, C529|Vagina|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C510-C512,C518, C529|Vagina|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C510-C512,C518, C529|Vagina|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C510-C512,C518, C529|Vagina|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C510-C512,C518, C529|Vagina|898|Carcinosarcoma|8980/3|Carcinosarcoma
C510-C512,C518, C529|Vagina|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C510-C512,C518, C529|Vagina|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C510-C512,C518, C529|Vagina|911|Mesonephroma|9110/3|Mesonephroma
C510-C512,C518, C529|Vagina|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C510-C512,C518, C529|Vagina|959|Lymphoma|9590/3|Lymphoma
C510-C512,C518, C529|Vagina|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C510-C512,C518, C529|Vagina|959|Lymphoma|9596/3|CompositeLymphoma
C510-C512,C518, C529|Vagina|959|Lymphoma|9597/3|CrostisDisease
C510-C512,C518, C529|Vagina|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C510-C512,C518, C529|Vagina|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C510-C512,C518, C529|Vagina|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C510-C512,C518, C529|Vagina|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C510-C512,C518, C529|Vagina|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C510-C512,C518, C529|Vagina|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C510-C512,C518, C529|Vagina|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C510-C512,C518, C529|Vagina|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C510-C512,C518, C529|Vagina|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C510-C512,C518, C529|Vagina|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C510-C512,C518, C529|Vagina|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C510-C512,C518, C529|Vagina|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C510-C512,C518, C529|Vagina|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C510-C512,C518, C529|Vagina|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C510-C512,C518, C529|Vagina|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C510-C512,C518, C529|Vagina|967|BCellLymphomas|9673/3|MantleCellLymphoma
C510-C512,C518, C529|Vagina|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C510-C512,C518, C529|Vagina|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C510-C512,C518, C529|Vagina|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C510-C512,C518, C529|Vagina|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C510-C512,C518, C529|Vagina|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C510-C512,C518, C529|Vagina|969|FollicularAdenoma|9690/3|LymphomaFollicular
C510-C512,C518, C529|Vagina|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C510-C512,C518, C529|Vagina|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C510-C512,C518, C529|Vagina|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C510-C512,C518, C529|Vagina|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C510-C512,C518, C529|Vagina|970|TCellLymphoma|9700/3|MycosisFungoides
C510-C512,C518, C529|Vagina|970|TCellLymphoma|9701/3|SezarySyndrome
C510-C512,C518, C529|Vagina|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C510-C512,C518, C529|Vagina|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C510-C512,C518, C529|Vagina|970|TCellLymphoma|9708/3|TCellLymphoma
C510-C512,C518, C529|Vagina|970|TCellLymphoma|9709/3|CutaneousTCellNonHodgkinLymphoma
C510-C512,C518, C529|Vagina|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C510-C512,C518, C529|Vagina|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C510-C512,C518, C529|Vagina|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C510-C512,C518, C529|Vagina|971|AdultNonHodgkinLymphoma|9718/3|CALCL
C510-C512,C518, C529|Vagina|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C510-C512,C518, C529|Vagina|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C510-C512,C518, C529|Vagina|972|LymphoblasticLymphoma|9725/3|HydroaVacciniformeLikeLymphoma
C510-C512,C518, C529|Vagina|972|LymphoblasticLymphoma|9726/3|TCellLymphoma
C510-C512,C518, C529|Vagina|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C510-C512,C518, C529|Vagina|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C510-C512,C518, C529|Vagina|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9731/3|Plasmacytoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C510-C512,C518, C529|Vagina|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C510-C512,C518, C529|Vagina|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C510-C512,C518, C529|Vagina|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C510-C512,C518, C529|Vagina|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C510-C512,C518, C529|Vagina|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C510-C512,C518, C529|Vagina|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C510-C512,C518, C529|Vagina|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C510-C512,C518, C529|Vagina|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C510-C512,C518, C529|Vagina|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C510-C512,C518, C529|Vagina|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C510-C512,C518, C529|Vagina|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C510-C512,C518, C529|Vagina|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9812/3|null
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9813/3|null
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9814/3|null
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9817/3|null
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9818/3|null
C510-C512,C518, C529|Vagina|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C510-C512,C518, C529|Vagina|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C510-C512,C518, C529|Vagina|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C510-C512,C518, C529|Vagina|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C510-C512,C518, C529|Vagina|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C510-C512,C518, C529|Vagina|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C510-C512,C518, C529|Vagina|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C510-C512,C518, C529|Vagina|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C519|Vulva|801|Carcinoma|8010/2|InSituCancer
C519|Vulva|801|Carcinoma|8010/3|CarcinomaNOSDNE
C519|Vulva|801|Carcinoma|8011/3|MalignantEpithelioma
C519|Vulva|801|Carcinoma|8012/3|LargeCellCarcinoma
C519|Vulva|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C519|Vulva|801|Carcinoma|8014/3|LargeCellCarcinoma
C519|Vulva|801|Carcinoma|8015/3|GlassyCellCarcinoma
C519|Vulva|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C519|Vulva|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C519|Vulva|802|Carcinoma|8022/3|PleomorphicCarcinoma
C519|Vulva|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C519|Vulva|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C519|Vulva|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C519|Vulva|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C519|Vulva|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C519|Vulva|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C519|Vulva|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8071/2|KeratinizingSquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C519|Vulva|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C519|Vulva|807|SquamousCellCarcinoma|8077/2|IntraepithelialNeoplasia
C519|Vulva|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C519|Vulva|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C519|Vulva|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C519|Vulva|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C519|Vulva|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C519|Vulva|809|BasalCellCarcinoma|8090/3|BasalCellCarcinoma
C519|Vulva|809|BasalCellCarcinoma|8091/3|SuperficialBasalCellCarcinoma
C519|Vulva|809|BasalCellCarcinoma|8092/3|SkinInfiltratingBasalCellCarcinoma
C519|Vulva|809|BasalCellCarcinoma|8093/3|FibroepitheliomaOfPinkus
C519|Vulva|809|BasalCellCarcinoma|8094/3|SkinBasosquamousCellCarcinoma
C519|Vulva|809|BasalCellCarcinoma|8095/3|SkinMetatypicalCarcinoma
C519|Vulva|809|BasalCellCarcinoma|8097/3|SkinNodularBasalCellCarcinoma
C519|Vulva|809|BasalCellCarcinoma|8098/3|SkinAdenoidBasalCellCarcinoma
C519|Vulva|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C519|Vulva|811|PilomatricalCarcinoma|8110/3|PilomatricalCarcinoma
C519|Vulva|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C519|Vulva|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C519|Vulva|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C519|Vulva|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C519|Vulva|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C519|Vulva|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C519|Vulva|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C519|Vulva|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C519|Vulva|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C519|Vulva|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C519|Vulva|814|Adenocarcinoma|8140/3|Adenocarcinoma
C519|Vulva|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C519|Vulva|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C519|Vulva|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C519|Vulva|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C519|Vulva|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C519|Vulva|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C519|Vulva|824|AtypicalCarcinoidTumor|8247/3|MerkelCellCarcinoma
C519|Vulva|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C519|Vulva|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C519|Vulva|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C519|Vulva|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C519|Vulva|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C519|Vulva|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C519|Vulva|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C519|Vulva|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C519|Vulva|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C519|Vulva|838|CarcinomaEndometrioid|8380/3|CarcinomaEndometrioid
C519|Vulva|839|AdnexalCarcinoma|8390/3|AdnexalCarcinoma
C519|Vulva|840|SweatGlandAdenocarcinoma|8400/3|SweatGlandAdenocarcinoma
C519|Vulva|840|SweatGlandAdenocarcinoma|8401/3|ApocrineAdenocarcinoma
C519|Vulva|841|EccrineAdenocarcinoma|8410/3|SebaceousAdenocarcinoma
C519|Vulva|841|EccrineAdenocarcinoma|8413/3|EccrineAdenocarcinoma
C519|Vulva|842|CeruminousAdenocarcinoma|8420/3|CeruminousAdenocarcinoma
C519|Vulva|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C519|Vulva|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C519|Vulva|848|MucinousAdenocarcinoma|8482/3|AdenocarcinomaEndocervicalType
C519|Vulva|854|PagetDiseaseExtramammary|8542/3|PagetDiseaseExtramammary
C519|Vulva|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C519|Vulva|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C519|Vulva|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C519|Vulva|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C519|Vulva|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C519|Vulva|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C519|Vulva|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C519|Vulva|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C519|Vulva|872|Melanoma|8720/2|Stage0SkinMelanoma
C519|Vulva|872|Melanoma|8720/3|Melanoma
C519|Vulva|872|Melanoma|8721/3|NodularMelanoma
C519|Vulva|872|Melanoma|8722/3|BalloonCellMelanoma
C519|Vulva|872|Melanoma|8723/3|RegressingMelanoma
C519|Vulva|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C519|Vulva|874|Nevus|8740/3|MelanomaInJunctionalNevus
C519|Vulva|874|Nevus|8741/2|PrecancerousMelanosis
C519|Vulva|874|Nevus|8741/3|Melanoma
C519|Vulva|874|Nevus|8742/2|LentigoMaligna
C519|Vulva|874|Nevus|8742/3|LentigoMalignaMelanoma
C519|Vulva|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C519|Vulva|874|Nevus|8745/3|DesmoplasticMelanoma
C519|Vulva|874|Nevus|8746/3|MucosalLentiginousMelanoma
C519|Vulva|876|Nevus|8761/3|GiantCongenitalNevus
C519|Vulva|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C519|Vulva|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C519|Vulva|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C519|Vulva|878|MelanomaArisingFromBlueNevus|8780/3|MelanomaArisingFromBlueNevus
C519|Vulva|880|Sarcoma|8800/3|Sarcoma
C519|Vulva|880|Sarcoma|8801/3|SpindleCellSarcoma
C519|Vulva|880|Sarcoma|8802/3|GiantCellSarcoma
C519|Vulva|880|Sarcoma|8803/3|SmallCellSarcoma
C519|Vulva|880|Sarcoma|8804/3|SarcomaEpithelioid
C519|Vulva|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C519|Vulva|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C519|Vulva|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C519|Vulva|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C519|Vulva|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C519|Vulva|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C519|Vulva|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C519|Vulva|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C519|Vulva|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C519|Vulva|883|BenignFibrousHistiocytoma|8832/3|DermatofibrosarcomaProtuberans
C519|Vulva|885|Liposarcoma|8850/3|Liposarcoma
C519|Vulva|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C519|Vulva|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C519|Vulva|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C519|Vulva|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C519|Vulva|885|Liposarcoma|8855/3|Liposarcoma
C519|Vulva|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C519|Vulva|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C519|Vulva|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C519|Vulva|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C519|Vulva|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C519|Vulva|889|MyomatousNeoplasm|8895/3|Myosarcoma
C519|Vulva|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C519|Vulva|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C519|Vulva|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C519|Vulva|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C519|Vulva|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C519|Vulva|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C519|Vulva|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C519|Vulva|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C519|Vulva|898|Carcinosarcoma|8980/3|Carcinosarcoma
C519|Vulva|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C519|Vulva|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C519|Vulva|911|Mesonephroma|9110/3|Mesonephroma
C519|Vulva|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C519|Vulva|959|Lymphoma|9590/3|Lymphoma
C519|Vulva|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C519|Vulva|959|Lymphoma|9596/3|CompositeLymphoma
C519|Vulva|959|Lymphoma|9597/3|CrostisDisease
C519|Vulva|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C519|Vulva|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C519|Vulva|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C519|Vulva|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C519|Vulva|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C519|Vulva|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C519|Vulva|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C519|Vulva|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C519|Vulva|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C519|Vulva|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C519|Vulva|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C519|Vulva|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C519|Vulva|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C519|Vulva|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C519|Vulva|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C519|Vulva|967|BCellLymphomas|9673/3|MantleCellLymphoma
C519|Vulva|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C519|Vulva|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C519|Vulva|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C519|Vulva|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C519|Vulva|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C519|Vulva|969|FollicularAdenoma|9690/3|LymphomaFollicular
C519|Vulva|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C519|Vulva|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C519|Vulva|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C519|Vulva|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C519|Vulva|970|TCellLymphoma|9700/3|MycosisFungoides
C519|Vulva|970|TCellLymphoma|9701/3|SezarySyndrome
C519|Vulva|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C519|Vulva|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C519|Vulva|970|TCellLymphoma|9708/3|TCellLymphoma
C519|Vulva|970|TCellLymphoma|9709/3|CutaneousTCellNonHodgkinLymphoma
C519|Vulva|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C519|Vulva|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C519|Vulva|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C519|Vulva|971|AdultNonHodgkinLymphoma|9718/3|CALCL
C519|Vulva|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C519|Vulva|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C519|Vulva|972|LymphoblasticLymphoma|9725/3|HydroaVacciniformeLikeLymphoma
C519|Vulva|972|LymphoblasticLymphoma|9726/3|TCellLymphoma
C519|Vulva|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C519|Vulva|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C519|Vulva|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C519|Vulva|973|Plasmacytoma|9731/3|Plasmacytoma
C519|Vulva|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C519|Vulva|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C519|Vulva|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C519|Vulva|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C519|Vulva|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C519|Vulva|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C519|Vulva|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C519|Vulva|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C519|Vulva|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C519|Vulva|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C519|Vulva|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C519|Vulva|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C519|Vulva|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C519|Vulva|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C519|Vulva|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C519|Vulva|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C519|Vulva|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C519|Vulva|981|PrecursorLymphoidNeoplasm|9812/3|null
C519|Vulva|981|PrecursorLymphoidNeoplasm|9813/3|null
C519|Vulva|981|PrecursorLymphoidNeoplasm|9814/3|null
C519|Vulva|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C519|Vulva|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C519|Vulva|981|PrecursorLymphoidNeoplasm|9817/3|null
C519|Vulva|981|PrecursorLymphoidNeoplasm|9818/3|null
C519|Vulva|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C519|Vulva|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C519|Vulva|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C519|Vulva|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C519|Vulva|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C519|Vulva|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C519|Vulva|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C519|Vulva|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C530-C531,C538-C539|CervixUteri|801|Carcinoma|8010/2|InSituCancer
C530-C531,C538-C539|CervixUteri|801|Carcinoma|8010/3|CarcinomaNOSDNE
C530-C531,C538-C539|CervixUteri|801|Carcinoma|8011/3|MalignantEpithelioma
C530-C531,C538-C539|CervixUteri|801|Carcinoma|8012/3|LargeCellCarcinoma
C530-C531,C538-C539|CervixUteri|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C530-C531,C538-C539|CervixUteri|801|Carcinoma|8014/3|LargeCellCarcinoma
C530-C531,C538-C539|CervixUteri|801|Carcinoma|8015/3|GlassyCellCarcinoma
C530-C531,C538-C539|CervixUteri|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C530-C531,C538-C539|CervixUteri|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C530-C531,C538-C539|CervixUteri|802|Carcinoma|8022/3|PleomorphicCarcinoma
C530-C531,C538-C539|CervixUteri|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C530-C531,C538-C539|CervixUteri|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C530-C531,C538-C539|CervixUteri|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C530-C531,C538-C539|CervixUteri|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C530-C531,C538-C539|CervixUteri|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C530-C531,C538-C539|CervixUteri|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C530-C531,C538-C539|CervixUteri|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C530-C531,C538-C539|CervixUteri|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C530-C531,C538-C539|CervixUteri|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C530-C531,C538-C539|CervixUteri|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C530-C531,C538-C539|CervixUteri|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C530-C531,C538-C539|CervixUteri|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C530-C531,C538-C539|CervixUteri|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8071/2|KeratinizingSquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8072/2|NonkeratinisingSquamousCellCarcinomaInSituDNE
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8077/2|IntraepithelialNeoplasia
C530-C531,C538-C539|CervixUteri|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C530-C531,C538-C539|CervixUteri|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C530-C531,C538-C539|CervixUteri|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C530-C531,C538-C539|CervixUteri|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C530-C531,C538-C539|CervixUteri|809|BasalCellCarcinoma|8098/3|SkinAdenoidBasalCellCarcinoma
C530-C531,C538-C539|CervixUteri|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C530-C531,C538-C539|CervixUteri|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C530-C531,C538-C539|CervixUteri|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C530-C531,C538-C539|CervixUteri|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C530-C531,C538-C539|CervixUteri|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C530-C531,C538-C539|CervixUteri|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C530-C531,C538-C539|CervixUteri|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C530-C531,C538-C539|CervixUteri|814|Adenocarcinoma|8140/3|Adenocarcinoma
C530-C531,C538-C539|CervixUteri|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C530-C531,C538-C539|CervixUteri|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C530-C531,C538-C539|CervixUteri|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C530-C531,C538-C539|CervixUteri|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C530-C531,C538-C539|CervixUteri|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C530-C531,C538-C539|CervixUteri|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C530-C531,C538-C539|CervixUteri|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C530-C531,C538-C539|CervixUteri|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C530-C531,C538-C539|CervixUteri|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C530-C531,C538-C539|CervixUteri|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C530-C531,C538-C539|CervixUteri|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C530-C531,C538-C539|CervixUteri|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C530-C531,C538-C539|CervixUteri|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C530-C531,C538-C539|CervixUteri|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C530-C531,C538-C539|CervixUteri|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C530-C531,C538-C539|CervixUteri|838|CarcinomaEndometrioid|8384/3|AdenocarcinomaEndocervicalType
C530-C531,C538-C539|CervixUteri|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C530-C531,C538-C539|CervixUteri|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C530-C531,C538-C539|CervixUteri|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C530-C531,C538-C539|CervixUteri|848|MucinousAdenocarcinoma|8482/3|AdenocarcinomaEndocervicalType
C530-C531,C538-C539|CervixUteri|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C530-C531,C538-C539|CervixUteri|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C530-C531,C538-C539|CervixUteri|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C530-C531,C538-C539|CervixUteri|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C530-C531,C538-C539|CervixUteri|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C530-C531,C538-C539|CervixUteri|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C530-C531,C538-C539|CervixUteri|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C530-C531,C538-C539|CervixUteri|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C530-C531,C538-C539|CervixUteri|880|Sarcoma|8800/3|Sarcoma
C530-C531,C538-C539|CervixUteri|880|Sarcoma|8801/3|SpindleCellSarcoma
C530-C531,C538-C539|CervixUteri|880|Sarcoma|8802/3|GiantCellSarcoma
C530-C531,C538-C539|CervixUteri|880|Sarcoma|8803/3|SmallCellSarcoma
C530-C531,C538-C539|CervixUteri|880|Sarcoma|8804/3|SarcomaEpithelioid
C530-C531,C538-C539|CervixUteri|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C530-C531,C538-C539|CervixUteri|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C530-C531,C538-C539|CervixUteri|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C530-C531,C538-C539|CervixUteri|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C530-C531,C538-C539|CervixUteri|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C530-C531,C538-C539|CervixUteri|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C530-C531,C538-C539|CervixUteri|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C530-C531,C538-C539|CervixUteri|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C530-C531,C538-C539|CervixUteri|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C530-C531,C538-C539|CervixUteri|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C530-C531,C538-C539|CervixUteri|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C530-C531,C538-C539|CervixUteri|889|MyomatousNeoplasm|8895/3|Myosarcoma
C530-C531,C538-C539|CervixUteri|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C530-C531,C538-C539|CervixUteri|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C530-C531,C538-C539|CervixUteri|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C530-C531,C538-C539|CervixUteri|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C530-C531,C538-C539|CervixUteri|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C530-C531,C538-C539|CervixUteri|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C530-C531,C538-C539|CervixUteri|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C530-C531,C538-C539|CervixUteri|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C530-C531,C538-C539|CervixUteri|898|Carcinosarcoma|8980/3|Carcinosarcoma
C530-C531,C538-C539|CervixUteri|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C530-C531,C538-C539|CervixUteri|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C530-C531,C538-C539|CervixUteri|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C530-C531,C538-C539|CervixUteri|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C530-C531,C538-C539|CervixUteri|911|Mesonephroma|9110/3|Mesonephroma
C530-C531,C538-C539|CervixUteri|959|Lymphoma|9590/3|Lymphoma
C530-C531,C538-C539|CervixUteri|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C530-C531,C538-C539|CervixUteri|959|Lymphoma|9596/3|CompositeLymphoma
C530-C531,C538-C539|CervixUteri|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C530-C531,C538-C539|CervixUteri|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C530-C531,C538-C539|CervixUteri|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C530-C531,C538-C539|CervixUteri|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C530-C531,C538-C539|CervixUteri|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C530-C531,C538-C539|CervixUteri|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C530-C531,C538-C539|CervixUteri|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C530-C531,C538-C539|CervixUteri|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C530-C531,C538-C539|CervixUteri|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C530-C531,C538-C539|CervixUteri|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C530-C531,C538-C539|CervixUteri|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C530-C531,C538-C539|CervixUteri|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C530-C531,C538-C539|CervixUteri|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C530-C531,C538-C539|CervixUteri|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C530-C531,C538-C539|CervixUteri|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C530-C531,C538-C539|CervixUteri|967|BCellLymphomas|9673/3|MantleCellLymphoma
C530-C531,C538-C539|CervixUteri|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C530-C531,C538-C539|CervixUteri|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C530-C531,C538-C539|CervixUteri|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C530-C531,C538-C539|CervixUteri|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C530-C531,C538-C539|CervixUteri|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C530-C531,C538-C539|CervixUteri|969|FollicularAdenoma|9690/3|LymphomaFollicular
C530-C531,C538-C539|CervixUteri|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C530-C531,C538-C539|CervixUteri|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C530-C531,C538-C539|CervixUteri|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C530-C531,C538-C539|CervixUteri|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C530-C531,C538-C539|CervixUteri|970|TCellLymphoma|9701/3|SezarySyndrome
C530-C531,C538-C539|CervixUteri|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C530-C531,C538-C539|CervixUteri|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C530-C531,C538-C539|CervixUteri|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C530-C531,C538-C539|CervixUteri|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C530-C531,C538-C539|CervixUteri|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C530-C531,C538-C539|CervixUteri|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C530-C531,C538-C539|CervixUteri|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C530-C531,C538-C539|CervixUteri|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C530-C531,C538-C539|CervixUteri|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C530-C531,C538-C539|CervixUteri|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C530-C531,C538-C539|CervixUteri|973|Plasmacytoma|9731/3|Plasmacytoma
C530-C531,C538-C539|CervixUteri|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C530-C531,C538-C539|CervixUteri|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C530-C531,C538-C539|CervixUteri|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C530-C531,C538-C539|CervixUteri|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C530-C531,C538-C539|CervixUteri|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C530-C531,C538-C539|CervixUteri|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C530-C531,C538-C539|CervixUteri|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C530-C531,C538-C539|CervixUteri|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C530-C531,C538-C539|CervixUteri|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C530-C531,C538-C539|CervixUteri|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C530-C531,C538-C539|CervixUteri|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C530-C531,C538-C539|CervixUteri|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C530-C531,C538-C539|CervixUteri|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C530-C531,C538-C539|CervixUteri|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C530-C531,C538-C539|CervixUteri|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C530-C531,C538-C539|CervixUteri|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9812/3|null
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9813/3|null
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9814/3|null
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9817/3|null
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9818/3|null
C530-C531,C538-C539|CervixUteri|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C530-C531,C538-C539|CervixUteri|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C530-C531,C538-C539|CervixUteri|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C530-C531,C538-C539|CervixUteri|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C530-C531,C538-C539|CervixUteri|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C530-C531,C538-C539|CervixUteri|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C530-C531,C538-C539|CervixUteri|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C530-C531,C538-C539|CervixUteri|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C540-C543,C548-C549|CorpusUteri|801|Carcinoma|8010/2|InSituCancer
C540-C543,C548-C549|CorpusUteri|801|Carcinoma|8010/3|CarcinomaNOSDNE
C540-C543,C548-C549|CorpusUteri|801|Carcinoma|8011/3|MalignantEpithelioma
C540-C543,C548-C549|CorpusUteri|801|Carcinoma|8012/3|LargeCellCarcinoma
C540-C543,C548-C549|CorpusUteri|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C540-C543,C548-C549|CorpusUteri|801|Carcinoma|8014/3|LargeCellCarcinoma
C540-C543,C548-C549|CorpusUteri|801|Carcinoma|8015/3|GlassyCellCarcinoma
C540-C543,C548-C549|CorpusUteri|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C540-C543,C548-C549|CorpusUteri|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C540-C543,C548-C549|CorpusUteri|802|Carcinoma|8022/3|PleomorphicCarcinoma
C540-C543,C548-C549|CorpusUteri|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C540-C543,C548-C549|CorpusUteri|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C540-C543,C548-C549|CorpusUteri|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C540-C543,C548-C549|CorpusUteri|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C540-C543,C548-C549|CorpusUteri|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C540-C543,C548-C549|CorpusUteri|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C540-C543,C548-C549|CorpusUteri|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C540-C543,C548-C549|CorpusUteri|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C540-C543,C548-C549|CorpusUteri|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C540-C543,C548-C549|CorpusUteri|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C540-C543,C548-C549|CorpusUteri|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C540-C543,C548-C549|CorpusUteri|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C540-C543,C548-C549|CorpusUteri|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C540-C543,C548-C549|CorpusUteri|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C540-C543,C548-C549|CorpusUteri|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C540-C543,C548-C549|CorpusUteri|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C540-C543,C548-C549|CorpusUteri|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C540-C543,C548-C549|CorpusUteri|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C540-C543,C548-C549|CorpusUteri|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C540-C543,C548-C549|CorpusUteri|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C540-C543,C548-C549|CorpusUteri|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C540-C543,C548-C549|CorpusUteri|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C540-C543,C548-C549|CorpusUteri|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C540-C543,C548-C549|CorpusUteri|814|Adenocarcinoma|8140/3|Adenocarcinoma
C540-C543,C548-C549|CorpusUteri|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C540-C543,C548-C549|CorpusUteri|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C540-C543,C548-C549|CorpusUteri|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C540-C543,C548-C549|CorpusUteri|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|823|SolidCarcinoma|8230/2|InSituCancer
C540-C543,C548-C549|CorpusUteri|823|SolidCarcinoma|8230/3|SolidCarcinoma
C540-C543,C548-C549|CorpusUteri|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C540-C543,C548-C549|CorpusUteri|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C540-C543,C548-C549|CorpusUteri|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C540-C543,C548-C549|CorpusUteri|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C540-C543,C548-C549|CorpusUteri|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C540-C543,C548-C549|CorpusUteri|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C540-C543,C548-C549|CorpusUteri|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C540-C543,C548-C549|CorpusUteri|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|838|CarcinomaEndometrioid|8380/2|AtypicalEndometrialHyperplasia
C540-C543,C548-C549|CorpusUteri|838|CarcinomaEndometrioid|8380/3|CarcinomaEndometrioid
C540-C543,C548-C549|CorpusUteri|838|CarcinomaEndometrioid|8381/3|EndometrioidAdenofibromaMalignant
C540-C543,C548-C549|CorpusUteri|838|CarcinomaEndometrioid|8382/3|CarcinomaEndometrioid
C540-C543,C548-C549|CorpusUteri|838|CarcinomaEndometrioid|8383/3|CarcinomaEndometrioid
C540-C543,C548-C549|CorpusUteri|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C540-C543,C548-C549|CorpusUteri|844|Cystadenocarcinoma|8441/1|SerousAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|844|Cystadenocarcinoma|8441/2|SerousTubalIntraepithelialCarcinoma
C540-C543,C548-C549|CorpusUteri|844|Cystadenocarcinoma|8441/3|SerousCystadenocarcinoma
C540-C543,C548-C549|CorpusUteri|846|PapillarySerousCystadenocarcinoma|8460/3|PapillarySerousCystadenocarcinoma
C540-C543,C548-C549|CorpusUteri|846|PapillarySerousCystadenocarcinoma|8461/3|SerousSurfacePapillaryCarcinoma
C540-C543,C548-C549|CorpusUteri|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|848|MucinousAdenocarcinoma|8482/3|AdenocarcinomaEndocervicalType
C540-C543,C548-C549|CorpusUteri|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C540-C543,C548-C549|CorpusUteri|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C540-C543,C548-C549|CorpusUteri|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C540-C543,C548-C549|CorpusUteri|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C540-C543,C548-C549|CorpusUteri|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C540-C543,C548-C549|CorpusUteri|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C540-C543,C548-C549|CorpusUteri|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C540-C543,C548-C549|CorpusUteri|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C540-C543,C548-C549|CorpusUteri|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C540-C543,C548-C549|CorpusUteri|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C540-C543,C548-C549|CorpusUteri|880|Sarcoma|8800/3|Sarcoma
C540-C543,C548-C549|CorpusUteri|880|Sarcoma|8801/3|SpindleCellSarcoma
C540-C543,C548-C549|CorpusUteri|880|Sarcoma|8802/3|GiantCellSarcoma
C540-C543,C548-C549|CorpusUteri|880|Sarcoma|8803/3|SmallCellSarcoma
C540-C543,C548-C549|CorpusUteri|880|Sarcoma|8804/3|SarcomaEpithelioid
C540-C543,C548-C549|CorpusUteri|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C540-C543,C548-C549|CorpusUteri|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C540-C543,C548-C549|CorpusUteri|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C540-C543,C548-C549|CorpusUteri|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C540-C543,C548-C549|CorpusUteri|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C540-C543,C548-C549|CorpusUteri|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C540-C543,C548-C549|CorpusUteri|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C540-C543,C548-C549|CorpusUteri|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C540-C543,C548-C549|CorpusUteri|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C540-C543,C548-C549|CorpusUteri|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C540-C543,C548-C549|CorpusUteri|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C540-C543,C548-C549|CorpusUteri|889|MyomatousNeoplasm|8895/3|Myosarcoma
C540-C543,C548-C549|CorpusUteri|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C540-C543,C548-C549|CorpusUteri|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C540-C543,C548-C549|CorpusUteri|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C540-C543,C548-C549|CorpusUteri|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C540-C543,C548-C549|CorpusUteri|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C540-C543,C548-C549|CorpusUteri|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C540-C543,C548-C549|CorpusUteri|893|StromalSarcoma|8930/3|EndometrialStromalSarcoma
C540-C543,C548-C549|CorpusUteri|893|StromalSarcoma|8931/3|LowGradeEndometrioidStromalSarcoma
C540-C543,C548-C549|CorpusUteri|893|StromalSarcoma|8933/3|Adenosarcoma
C540-C543,C548-C549|CorpusUteri|893|StromalSarcoma|8934/3|Carcinofibroma
C540-C543,C548-C549|CorpusUteri|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C540-C543,C548-C549|CorpusUteri|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C540-C543,C548-C549|CorpusUteri|898|Carcinosarcoma|8980/3|Carcinosarcoma
C540-C543,C548-C549|CorpusUteri|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C540-C543,C548-C549|CorpusUteri|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C540-C543,C548-C549|CorpusUteri|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C540-C543,C548-C549|CorpusUteri|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C540-C543,C548-C549|CorpusUteri|911|Mesonephroma|9110/3|Mesonephroma
C540-C543,C548-C549|CorpusUteri|959|Lymphoma|9590/3|Lymphoma
C540-C543,C548-C549|CorpusUteri|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C540-C543,C548-C549|CorpusUteri|959|Lymphoma|9596/3|CompositeLymphoma
C540-C543,C548-C549|CorpusUteri|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C540-C543,C548-C549|CorpusUteri|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C540-C543,C548-C549|CorpusUteri|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C540-C543,C548-C549|CorpusUteri|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C540-C543,C548-C549|CorpusUteri|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C540-C543,C548-C549|CorpusUteri|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C540-C543,C548-C549|CorpusUteri|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C540-C543,C548-C549|CorpusUteri|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C540-C543,C548-C549|CorpusUteri|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C540-C543,C548-C549|CorpusUteri|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C540-C543,C548-C549|CorpusUteri|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C540-C543,C548-C549|CorpusUteri|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C540-C543,C548-C549|CorpusUteri|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C540-C543,C548-C549|CorpusUteri|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C540-C543,C548-C549|CorpusUteri|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C540-C543,C548-C549|CorpusUteri|967|BCellLymphomas|9673/3|MantleCellLymphoma
C540-C543,C548-C549|CorpusUteri|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C540-C543,C548-C549|CorpusUteri|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C540-C543,C548-C549|CorpusUteri|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C540-C543,C548-C549|CorpusUteri|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C540-C543,C548-C549|CorpusUteri|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C540-C543,C548-C549|CorpusUteri|969|FollicularAdenoma|9690/3|LymphomaFollicular
C540-C543,C548-C549|CorpusUteri|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C540-C543,C548-C549|CorpusUteri|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C540-C543,C548-C549|CorpusUteri|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C540-C543,C548-C549|CorpusUteri|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C540-C543,C548-C549|CorpusUteri|970|TCellLymphoma|9701/3|SezarySyndrome
C540-C543,C548-C549|CorpusUteri|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C540-C543,C548-C549|CorpusUteri|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C540-C543,C548-C549|CorpusUteri|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C540-C543,C548-C549|CorpusUteri|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C540-C543,C548-C549|CorpusUteri|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C540-C543,C548-C549|CorpusUteri|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C540-C543,C548-C549|CorpusUteri|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C540-C543,C548-C549|CorpusUteri|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C540-C543,C548-C549|CorpusUteri|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C540-C543,C548-C549|CorpusUteri|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C540-C543,C548-C549|CorpusUteri|973|Plasmacytoma|9731/3|Plasmacytoma
C540-C543,C548-C549|CorpusUteri|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C540-C543,C548-C549|CorpusUteri|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C540-C543,C548-C549|CorpusUteri|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C540-C543,C548-C549|CorpusUteri|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C540-C543,C548-C549|CorpusUteri|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C540-C543,C548-C549|CorpusUteri|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C540-C543,C548-C549|CorpusUteri|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C540-C543,C548-C549|CorpusUteri|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C540-C543,C548-C549|CorpusUteri|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C540-C543,C548-C549|CorpusUteri|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C540-C543,C548-C549|CorpusUteri|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C540-C543,C548-C549|CorpusUteri|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C540-C543,C548-C549|CorpusUteri|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9812/3|null
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9813/3|null
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9814/3|null
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9817/3|null
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9818/3|null
C540-C543,C548-C549|CorpusUteri|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C540-C543,C548-C549|CorpusUteri|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C540-C543,C548-C549|CorpusUteri|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C540-C543,C548-C549|CorpusUteri|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C540-C543,C548-C549|CorpusUteri|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C540-C543,C548-C549|CorpusUteri|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C540-C543,C548-C549|CorpusUteri|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C540-C543,C548-C549|CorpusUteri|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C559|Uterus|801|Carcinoma|8010/2|InSituCancer
C559|Uterus|801|Carcinoma|8010/3|CarcinomaNOSDNE
C559|Uterus|801|Carcinoma|8011/3|MalignantEpithelioma
C559|Uterus|801|Carcinoma|8012/3|LargeCellCarcinoma
C559|Uterus|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C559|Uterus|801|Carcinoma|8014/3|LargeCellCarcinoma
C559|Uterus|801|Carcinoma|8015/3|GlassyCellCarcinoma
C559|Uterus|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C559|Uterus|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C559|Uterus|802|Carcinoma|8022/3|PleomorphicCarcinoma
C559|Uterus|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C559|Uterus|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C559|Uterus|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C559|Uterus|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C559|Uterus|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C559|Uterus|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C559|Uterus|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C559|Uterus|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C559|Uterus|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C559|Uterus|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C559|Uterus|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C559|Uterus|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C559|Uterus|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C559|Uterus|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C559|Uterus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C559|Uterus|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C559|Uterus|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C559|Uterus|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C559|Uterus|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C559|Uterus|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C559|Uterus|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C559|Uterus|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C559|Uterus|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C559|Uterus|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C559|Uterus|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C559|Uterus|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C559|Uterus|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C559|Uterus|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C559|Uterus|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C559|Uterus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C559|Uterus|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C559|Uterus|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C559|Uterus|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C559|Uterus|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C559|Uterus|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C559|Uterus|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C559|Uterus|821|AdenocarcinomaInAdenomatousPolyp|8210/2|AdenocarcinomaInSitu
C559|Uterus|821|AdenocarcinomaInAdenomatousPolyp|8210/3|AdenocarcinomaInAdenomatousPolyp
C559|Uterus|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C559|Uterus|823|SolidCarcinoma|8230/2|InSituCancer
C559|Uterus|823|SolidCarcinoma|8230/3|SolidCarcinoma
C559|Uterus|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C559|Uterus|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C559|Uterus|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C559|Uterus|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C559|Uterus|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C559|Uterus|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C559|Uterus|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C559|Uterus|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C559|Uterus|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C559|Uterus|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C559|Uterus|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C559|Uterus|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C559|Uterus|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C559|Uterus|844|Cystadenocarcinoma|8441/1|SerousAdenocarcinoma
C559|Uterus|844|Cystadenocarcinoma|8441/2|SerousTubalIntraepithelialCarcinoma
C559|Uterus|844|Cystadenocarcinoma|8441/3|SerousCystadenocarcinoma
C559|Uterus|846|PapillarySerousCystadenocarcinoma|8460/3|PapillarySerousCystadenocarcinoma
C559|Uterus|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C559|Uterus|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C559|Uterus|848|MucinousAdenocarcinoma|8482/3|AdenocarcinomaEndocervicalType
C559|Uterus|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C559|Uterus|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C559|Uterus|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C559|Uterus|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C559|Uterus|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C559|Uterus|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C559|Uterus|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C559|Uterus|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C559|Uterus|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C559|Uterus|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C559|Uterus|880|Sarcoma|8800/3|Sarcoma
C559|Uterus|880|Sarcoma|8801/3|SpindleCellSarcoma
C559|Uterus|880|Sarcoma|8802/3|GiantCellSarcoma
C559|Uterus|880|Sarcoma|8803/3|SmallCellSarcoma
C559|Uterus|880|Sarcoma|8804/3|SarcomaEpithelioid
C559|Uterus|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C559|Uterus|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C559|Uterus|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C559|Uterus|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C559|Uterus|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C559|Uterus|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C559|Uterus|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C559|Uterus|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C559|Uterus|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C559|Uterus|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C559|Uterus|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C559|Uterus|889|MyomatousNeoplasm|8895/3|Myosarcoma
C559|Uterus|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C559|Uterus|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C559|Uterus|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C559|Uterus|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C559|Uterus|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C559|Uterus|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C559|Uterus|893|StromalSarcoma|8930/3|EndometrialStromalSarcoma
C559|Uterus|893|StromalSarcoma|8931/3|LowGradeEndometrioidStromalSarcoma
C559|Uterus|893|StromalSarcoma|8934/3|Carcinofibroma
C559|Uterus|893|StromalSarcoma|8935/3|StromalSarcoma
C559|Uterus|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C559|Uterus|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C559|Uterus|898|Carcinosarcoma|8980/3|Carcinosarcoma
C559|Uterus|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C559|Uterus|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C559|Uterus|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C559|Uterus|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C559|Uterus|911|Mesonephroma|9110/3|Mesonephroma
C559|Uterus|959|Lymphoma|9590/3|Lymphoma
C559|Uterus|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C559|Uterus|959|Lymphoma|9596/3|CompositeLymphoma
C559|Uterus|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C559|Uterus|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C559|Uterus|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C559|Uterus|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C559|Uterus|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C559|Uterus|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C559|Uterus|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C559|Uterus|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C559|Uterus|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C559|Uterus|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C559|Uterus|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C559|Uterus|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C559|Uterus|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C559|Uterus|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C559|Uterus|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C559|Uterus|967|BCellLymphomas|9673/3|MantleCellLymphoma
C559|Uterus|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C559|Uterus|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C559|Uterus|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C559|Uterus|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C559|Uterus|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C559|Uterus|969|FollicularAdenoma|9690/3|LymphomaFollicular
C559|Uterus|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C559|Uterus|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C559|Uterus|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C559|Uterus|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C559|Uterus|970|TCellLymphoma|9701/3|SezarySyndrome
C559|Uterus|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C559|Uterus|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C559|Uterus|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C559|Uterus|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C559|Uterus|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C559|Uterus|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C559|Uterus|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C559|Uterus|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C559|Uterus|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C559|Uterus|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C559|Uterus|973|Plasmacytoma|9731/3|Plasmacytoma
C559|Uterus|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C559|Uterus|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C559|Uterus|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C559|Uterus|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C559|Uterus|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C559|Uterus|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C559|Uterus|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C559|Uterus|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C559|Uterus|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C559|Uterus|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C559|Uterus|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C559|Uterus|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C559|Uterus|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C559|Uterus|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C559|Uterus|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C559|Uterus|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C559|Uterus|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C559|Uterus|981|PrecursorLymphoidNeoplasm|9812/3|null
C559|Uterus|981|PrecursorLymphoidNeoplasm|9813/3|null
C559|Uterus|981|PrecursorLymphoidNeoplasm|9814/3|null
C559|Uterus|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C559|Uterus|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C559|Uterus|981|PrecursorLymphoidNeoplasm|9817/3|null
C559|Uterus|981|PrecursorLymphoidNeoplasm|9818/3|null
C559|Uterus|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C559|Uterus|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C559|Uterus|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C559|Uterus|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C559|Uterus|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C559|Uterus|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C559|Uterus|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C559|Uterus|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C569|Ovary|801|Carcinoma|8010/2|InSituCancer
C569|Ovary|801|Carcinoma|8010/3|CarcinomaNOSDNE
C569|Ovary|801|Carcinoma|8011/3|MalignantEpithelioma
C569|Ovary|801|Carcinoma|8012/3|LargeCellCarcinoma
C569|Ovary|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C569|Ovary|801|Carcinoma|8014/3|LargeCellCarcinoma
C569|Ovary|801|Carcinoma|8015/3|GlassyCellCarcinoma
C569|Ovary|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C569|Ovary|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C569|Ovary|802|Carcinoma|8022/3|PleomorphicCarcinoma
C569|Ovary|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C569|Ovary|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C569|Ovary|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C569|Ovary|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C569|Ovary|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C569|Ovary|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C569|Ovary|804|SmallCellCarcinoma|8041/3|OvarianSmallCellCarcinoma
C569|Ovary|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C569|Ovary|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C569|Ovary|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C569|Ovary|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C569|Ovary|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C569|Ovary|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C569|Ovary|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C569|Ovary|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C569|Ovary|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C569|Ovary|814|Adenocarcinoma|8140/3|Adenocarcinoma
C569|Ovary|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C569|Ovary|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C569|Ovary|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C569|Ovary|823|SolidCarcinoma|8230/2|InSituCancer
C569|Ovary|823|SolidCarcinoma|8230/3|SolidCarcinoma
C569|Ovary|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C569|Ovary|824|AtypicalCarcinoidTumor|8240/2|OvarianCarcinoidTumor
C569|Ovary|824|AtypicalCarcinoidTumor|8240/3|AtypicalCarcinoidTumor
C569|Ovary|824|AtypicalCarcinoidTumor|8241/3|ECCellCarcinoid
C569|Ovary|824|AtypicalCarcinoidTumor|8242/3|EnterochromaffinlikeCellCarcinoid
C569|Ovary|824|AtypicalCarcinoidTumor|8243/3|GobletCellCarcinoid
C569|Ovary|824|AtypicalCarcinoidTumor|8244/3|AdenocarcinoidTumor
C569|Ovary|824|AtypicalCarcinoidTumor|8245/3|AdenocarcinoidTumor
C569|Ovary|824|AtypicalCarcinoidTumor|8246/3|NeuroendocrineNeoplasm
C569|Ovary|824|AtypicalCarcinoidTumor|8249/3|AtypicalCarcinoidTumor
C569|Ovary|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C569|Ovary|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C569|Ovary|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C569|Ovary|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C569|Ovary|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C569|Ovary|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C569|Ovary|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C569|Ovary|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C569|Ovary|831|ClearCellAdenocarcinoma|8313/3|ClearCellAdenocarcinofibroma
C569|Ovary|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C569|Ovary|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C569|Ovary|838|CarcinomaEndometrioid|8380/3|CarcinomaEndometrioid
C569|Ovary|838|CarcinomaEndometrioid|8381/3|EndometrioidAdenofibromaMalignant
C569|Ovary|838|CarcinomaEndometrioid|8382/3|CarcinomaEndometrioid
C569|Ovary|838|CarcinomaEndometrioid|8383/3|CarcinomaEndometrioid
C569|Ovary|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C569|Ovary|844|Cystadenocarcinoma|8441/1|OvarianSerousCystadenocarcinoma
C569|Ovary|844|Cystadenocarcinoma|8441/2|SerousTubalIntraepithelialCarcinoma
C569|Ovary|844|Cystadenocarcinoma|8441/3|SerousCystadenocarcinoma
C569|Ovary|844|Cystadenocarcinoma|8442/1|SerousCystadenoma
C569|Ovary|845|PapillaryCystadenocarcinoma|8450/3|PapillaryCystadenocarcinoma
C569|Ovary|845|PapillaryCystadenocarcinoma|8451/1|PapillaryCystadenoma
C569|Ovary|846|PapillarySerousCystadenocarcinoma|8460/1|SerousAdenocarcinoma
C569|Ovary|846|PapillarySerousCystadenocarcinoma|8460/2|SerousCystadenocarcinoma
C569|Ovary|846|PapillarySerousCystadenocarcinoma|8460/3|PapillarySerousCystadenocarcinoma
C569|Ovary|846|PapillarySerousCystadenocarcinoma|8461/3|SerousSurfacePapillaryCarcinoma
C569|Ovary|846|PapillarySerousCystadenocarcinoma|8462/1|PapillaryCysticNeoplasm
C569|Ovary|847|MucinousCystadenocarcinoma|8470/2|MucinousCystadenocarcinoma
C569|Ovary|847|MucinousCystadenocarcinoma|8470/3|MucinousCystadenocarcinoma
C569|Ovary|847|MucinousCystadenocarcinoma|8471/3|PapillaryMucinousCystadenocarcinoma
C569|Ovary|847|MucinousCystadenocarcinoma|8472/1|CysticNeoplasm
C569|Ovary|847|MucinousCystadenocarcinoma|8473/1|PapillaryMucinousCystadenoma
C569|Ovary|847|MucinousCystadenocarcinoma|8474/3|OvarianSeromucinousTumor
C569|Ovary|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C569|Ovary|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C569|Ovary|848|MucinousAdenocarcinoma|8482/3|AdenocarcinomaEndocervicalType
C569|Ovary|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C569|Ovary|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C569|Ovary|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C569|Ovary|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C569|Ovary|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C569|Ovary|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C569|Ovary|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C569|Ovary|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C569|Ovary|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C569|Ovary|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C569|Ovary|859|OvarianSexCordStromalTumor|8590/3|OvarianSexCordStromalTumor
C569|Ovary|860|MalignantOvarianThecoma|8600/3|MalignantOvarianThecoma
C569|Ovary|862|GranulosaCellTumor|8620/3|MalignantGranulosaCellTumor
C569|Ovary|862|GranulosaCellTumor|8621/3|GranulosaCellThecaCellTumor
C569|Ovary|863|GonadalNeoplasm|8630/3|MalignantSertoliCellTumor
C569|Ovary|863|GonadalNeoplasm|8631/3|SertoliLeydigCellTumor
C569|Ovary|863|GonadalNeoplasm|8632/3|OvarianGynandroblastoma
C569|Ovary|863|GonadalNeoplasm|8634/3|SertoliLeydigCellTumor
C569|Ovary|867|SteroidCellTumorMalignant|8670/3|SteroidCellTumorMalignant
C569|Ovary|880|Sarcoma|8800/3|Sarcoma
C569|Ovary|880|Sarcoma|8801/3|SpindleCellSarcoma
C569|Ovary|880|Sarcoma|8802/3|GiantCellSarcoma
C569|Ovary|880|Sarcoma|8803/3|SmallCellSarcoma
C569|Ovary|880|Sarcoma|8804/3|SarcomaEpithelioid
C569|Ovary|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C569|Ovary|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C569|Ovary|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C569|Ovary|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C569|Ovary|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C569|Ovary|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C569|Ovary|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C569|Ovary|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C569|Ovary|884|Myxosarcoma|8840/3|Myxosarcoma
C569|Ovary|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C569|Ovary|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C569|Ovary|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C569|Ovary|889|MyomatousNeoplasm|8895/3|Myosarcoma
C569|Ovary|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C569|Ovary|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C569|Ovary|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C569|Ovary|898|Carcinosarcoma|8980/3|Carcinosarcoma
C569|Ovary|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C569|Ovary|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C569|Ovary|900|MalignantOvarianBrennerTumor|9000/3|MalignantOvarianBrennerTumor
C569|Ovary|901|Adenocarcinofibroma|9014/3|SerousAdenocarcinofibroma
C569|Ovary|901|Adenocarcinofibroma|9015/3|MucinousAdenocarcinofibroma
C569|Ovary|906|GermCellTumor|9060/3|Dysgerminoma
C569|Ovary|906|GermCellTumor|9064/3|Germinoma
C569|Ovary|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C569|Ovary|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C569|Ovary|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C569|Ovary|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C569|Ovary|908|Teratoma|9080/3|ImmatureTeratoma
C569|Ovary|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C569|Ovary|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C569|Ovary|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C569|Ovary|908|Teratoma|9084/3|Teratoma
C569|Ovary|908|Teratoma|9085/3|MixedGermCellTumor
C569|Ovary|909|MalignantStrumaOvarii|9090/3|MalignantStrumaOvarii
C569|Ovary|910|Choriocarcinoma|9100/3|Choriocarcinoma
C569|Ovary|910|Choriocarcinoma|9101/3|Choriocarcinoma
C569|Ovary|910|Choriocarcinoma|9105/3|EpithelioidTrophoblasticTumor
C569|Ovary|911|Mesonephroma|9110/3|Mesonephroma
C569|Ovary|959|Lymphoma|9590/3|Lymphoma
C569|Ovary|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C569|Ovary|959|Lymphoma|9596/3|CompositeLymphoma
C569|Ovary|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C569|Ovary|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C569|Ovary|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C569|Ovary|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C569|Ovary|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C569|Ovary|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C569|Ovary|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C569|Ovary|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C569|Ovary|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C569|Ovary|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C569|Ovary|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C569|Ovary|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C569|Ovary|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C569|Ovary|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C569|Ovary|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C569|Ovary|967|BCellLymphomas|9673/3|MantleCellLymphoma
C569|Ovary|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C569|Ovary|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C569|Ovary|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C569|Ovary|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C569|Ovary|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C569|Ovary|969|FollicularAdenoma|9690/3|LymphomaFollicular
C569|Ovary|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C569|Ovary|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C569|Ovary|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C569|Ovary|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C569|Ovary|970|TCellLymphoma|9701/3|SezarySyndrome
C569|Ovary|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C569|Ovary|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C569|Ovary|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C569|Ovary|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C569|Ovary|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C569|Ovary|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C569|Ovary|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C569|Ovary|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C569|Ovary|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C569|Ovary|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C569|Ovary|973|Plasmacytoma|9731/3|Plasmacytoma
C569|Ovary|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C569|Ovary|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C569|Ovary|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C569|Ovary|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C569|Ovary|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C569|Ovary|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C569|Ovary|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C569|Ovary|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C569|Ovary|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C569|Ovary|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C569|Ovary|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C569|Ovary|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C569|Ovary|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C569|Ovary|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C569|Ovary|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C569|Ovary|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C569|Ovary|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C569|Ovary|981|PrecursorLymphoidNeoplasm|9812/3|null
C569|Ovary|981|PrecursorLymphoidNeoplasm|9813/3|null
C569|Ovary|981|PrecursorLymphoidNeoplasm|9814/3|null
C569|Ovary|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C569|Ovary|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C569|Ovary|981|PrecursorLymphoidNeoplasm|9817/3|null
C569|Ovary|981|PrecursorLymphoidNeoplasm|9818/3|null
C569|Ovary|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C569|Ovary|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C569|Ovary|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C569|Ovary|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C569|Ovary|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C569|Ovary|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C569|Ovary|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C569|Ovary|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C570|FallopianTube|801|Carcinoma|8010/2|InSituCancer
C570|FallopianTube|801|Carcinoma|8010/3|CarcinomaNOSDNE
C570|FallopianTube|801|Carcinoma|8011/3|MalignantEpithelioma
C570|FallopianTube|801|Carcinoma|8012/3|LargeCellCarcinoma
C570|FallopianTube|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C570|FallopianTube|801|Carcinoma|8014/3|LargeCellCarcinoma
C570|FallopianTube|801|Carcinoma|8015/3|GlassyCellCarcinoma
C570|FallopianTube|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C570|FallopianTube|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C570|FallopianTube|802|Carcinoma|8022/3|PleomorphicCarcinoma
C570|FallopianTube|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C570|FallopianTube|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C570|FallopianTube|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C570|FallopianTube|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C570|FallopianTube|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C570|FallopianTube|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C570|FallopianTube|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C570|FallopianTube|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C570|FallopianTube|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C570|FallopianTube|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C570|FallopianTube|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C570|FallopianTube|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C570|FallopianTube|814|Adenocarcinoma|8140/3|Adenocarcinoma
C570|FallopianTube|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C570|FallopianTube|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C570|FallopianTube|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C570|FallopianTube|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C570|FallopianTube|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C570|FallopianTube|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C570|FallopianTube|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C570|FallopianTube|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C570|FallopianTube|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C570|FallopianTube|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C570|FallopianTube|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C570|FallopianTube|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C570|FallopianTube|838|CarcinomaEndometrioid|8380/3|CarcinomaEndometrioid
C570|FallopianTube|838|CarcinomaEndometrioid|8382/3|CarcinomaEndometrioid
C570|FallopianTube|838|CarcinomaEndometrioid|8383/3|CarcinomaEndometrioid
C570|FallopianTube|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C570|FallopianTube|844|Cystadenocarcinoma|8441/1|SerousAdenocarcinoma
C570|FallopianTube|844|Cystadenocarcinoma|8441/2|SerousTubalIntraepithelialCarcinoma
C570|FallopianTube|844|Cystadenocarcinoma|8441/3|SerousCystadenocarcinoma
C570|FallopianTube|846|PapillarySerousCystadenocarcinoma|8460/3|PapillarySerousCystadenocarcinoma
C570|FallopianTube|846|PapillarySerousCystadenocarcinoma|8461/3|SerousSurfacePapillaryCarcinoma
C570|FallopianTube|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C570|FallopianTube|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C570|FallopianTube|848|MucinousAdenocarcinoma|8482/3|AdenocarcinomaEndocervicalType
C570|FallopianTube|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C570|FallopianTube|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C570|FallopianTube|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C570|FallopianTube|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C570|FallopianTube|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C570|FallopianTube|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C570|FallopianTube|880|Sarcoma|8800/3|Sarcoma
C570|FallopianTube|880|Sarcoma|8801/3|SpindleCellSarcoma
C570|FallopianTube|880|Sarcoma|8802/3|GiantCellSarcoma
C570|FallopianTube|880|Sarcoma|8803/3|SmallCellSarcoma
C570|FallopianTube|880|Sarcoma|8804/3|SarcomaEpithelioid
C570|FallopianTube|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C570|FallopianTube|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C570|FallopianTube|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C570|FallopianTube|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C570|FallopianTube|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C570|FallopianTube|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C570|FallopianTube|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C570|FallopianTube|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C570|FallopianTube|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C570|FallopianTube|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C570|FallopianTube|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C570|FallopianTube|889|MyomatousNeoplasm|8895/3|Myosarcoma
C570|FallopianTube|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C570|FallopianTube|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C570|FallopianTube|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C570|FallopianTube|898|Carcinosarcoma|8980/3|Carcinosarcoma
C570|FallopianTube|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C570|FallopianTube|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C570|FallopianTube|911|Mesonephroma|9110/3|Mesonephroma
C570|FallopianTube|959|Lymphoma|9590/3|Lymphoma
C570|FallopianTube|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C570|FallopianTube|959|Lymphoma|9596/3|CompositeLymphoma
C570|FallopianTube|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C570|FallopianTube|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C570|FallopianTube|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C570|FallopianTube|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C570|FallopianTube|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C570|FallopianTube|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C570|FallopianTube|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C570|FallopianTube|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C570|FallopianTube|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C570|FallopianTube|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C570|FallopianTube|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C570|FallopianTube|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C570|FallopianTube|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C570|FallopianTube|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C570|FallopianTube|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C570|FallopianTube|967|BCellLymphomas|9673/3|MantleCellLymphoma
C570|FallopianTube|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C570|FallopianTube|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C570|FallopianTube|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C570|FallopianTube|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C570|FallopianTube|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C570|FallopianTube|969|FollicularAdenoma|9690/3|LymphomaFollicular
C570|FallopianTube|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C570|FallopianTube|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C570|FallopianTube|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C570|FallopianTube|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C570|FallopianTube|970|TCellLymphoma|9701/3|SezarySyndrome
C570|FallopianTube|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C570|FallopianTube|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C570|FallopianTube|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C570|FallopianTube|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C570|FallopianTube|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C570|FallopianTube|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C570|FallopianTube|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C570|FallopianTube|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C570|FallopianTube|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C570|FallopianTube|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C570|FallopianTube|973|Plasmacytoma|9731/3|Plasmacytoma
C570|FallopianTube|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C570|FallopianTube|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C570|FallopianTube|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C570|FallopianTube|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C570|FallopianTube|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C570|FallopianTube|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C570|FallopianTube|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C570|FallopianTube|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C570|FallopianTube|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C570|FallopianTube|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C570|FallopianTube|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C570|FallopianTube|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C570|FallopianTube|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C570|FallopianTube|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C570|FallopianTube|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C570|FallopianTube|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9812/3|null
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9813/3|null
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9814/3|null
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9817/3|null
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9818/3|null
C570|FallopianTube|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C570|FallopianTube|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C570|FallopianTube|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C570|FallopianTube|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C570|FallopianTube|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C570|FallopianTube|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C570|FallopianTube|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C570|FallopianTube|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C571-C574,C577-C579|FallopianTube|801|Carcinoma|8010/2|InSituCancer
C571-C574,C577-C579|FallopianTube|801|Carcinoma|8010/3|CarcinomaNOSDNE
C571-C574,C577-C579|FallopianTube|801|Carcinoma|8011/3|MalignantEpithelioma
C571-C574,C577-C579|FallopianTube|801|Carcinoma|8012/3|LargeCellCarcinoma
C571-C574,C577-C579|FallopianTube|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C571-C574,C577-C579|FallopianTube|801|Carcinoma|8014/3|LargeCellCarcinoma
C571-C574,C577-C579|FallopianTube|801|Carcinoma|8015/3|GlassyCellCarcinoma
C571-C574,C577-C579|FallopianTube|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C571-C574,C577-C579|FallopianTube|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C571-C574,C577-C579|FallopianTube|802|Carcinoma|8022/3|PleomorphicCarcinoma
C571-C574,C577-C579|FallopianTube|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C571-C574,C577-C579|FallopianTube|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C571-C574,C577-C579|FallopianTube|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C571-C574,C577-C579|FallopianTube|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C571-C574,C577-C579|FallopianTube|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C571-C574,C577-C579|FallopianTube|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C571-C574,C577-C579|FallopianTube|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C571-C574,C577-C579|FallopianTube|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C571-C574,C577-C579|FallopianTube|814|Adenocarcinoma|8140/3|Adenocarcinoma
C571-C574,C577-C579|FallopianTube|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C571-C574,C577-C579|FallopianTube|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C571-C574,C577-C579|FallopianTube|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C571-C574,C577-C579|FallopianTube|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C571-C574,C577-C579|FallopianTube|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C571-C574,C577-C579|FallopianTube|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C571-C574,C577-C579|FallopianTube|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C571-C574,C577-C579|FallopianTube|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C571-C574,C577-C579|FallopianTube|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C571-C574,C577-C579|FallopianTube|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C571-C574,C577-C579|FallopianTube|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C571-C574,C577-C579|FallopianTube|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C571-C574,C577-C579|FallopianTube|838|CarcinomaEndometrioid|8380/3|CarcinomaEndometrioid
C571-C574,C577-C579|FallopianTube|838|CarcinomaEndometrioid|8382/3|CarcinomaEndometrioid
C571-C574,C577-C579|FallopianTube|838|CarcinomaEndometrioid|8383/3|CarcinomaEndometrioid
C571-C574,C577-C579|FallopianTube|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C571-C574,C577-C579|FallopianTube|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C571-C574,C577-C579|FallopianTube|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C571-C574,C577-C579|FallopianTube|848|MucinousAdenocarcinoma|8482/3|AdenocarcinomaEndocervicalType
C571-C574,C577-C579|FallopianTube|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C571-C574,C577-C579|FallopianTube|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C571-C574,C577-C579|FallopianTube|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C571-C574,C577-C579|FallopianTube|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C571-C574,C577-C579|FallopianTube|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C571-C574,C577-C579|FallopianTube|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C571-C574,C577-C579|FallopianTube|880|Sarcoma|8800/3|Sarcoma
C571-C574,C577-C579|FallopianTube|880|Sarcoma|8801/3|SpindleCellSarcoma
C571-C574,C577-C579|FallopianTube|880|Sarcoma|8802/3|GiantCellSarcoma
C571-C574,C577-C579|FallopianTube|880|Sarcoma|8803/3|SmallCellSarcoma
C571-C574,C577-C579|FallopianTube|880|Sarcoma|8804/3|SarcomaEpithelioid
C571-C574,C577-C579|FallopianTube|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C571-C574,C577-C579|FallopianTube|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C571-C574,C577-C579|FallopianTube|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C571-C574,C577-C579|FallopianTube|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C571-C574,C577-C579|FallopianTube|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C571-C574,C577-C579|FallopianTube|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C571-C574,C577-C579|FallopianTube|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C571-C574,C577-C579|FallopianTube|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C571-C574,C577-C579|FallopianTube|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C571-C574,C577-C579|FallopianTube|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C571-C574,C577-C579|FallopianTube|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C571-C574,C577-C579|FallopianTube|889|MyomatousNeoplasm|8895/3|Myosarcoma
C571-C574,C577-C579|FallopianTube|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C571-C574,C577-C579|FallopianTube|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C571-C574,C577-C579|FallopianTube|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C571-C574,C577-C579|FallopianTube|898|Carcinosarcoma|8980/3|Carcinosarcoma
C571-C574,C577-C579|FallopianTube|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C571-C574,C577-C579|FallopianTube|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C571-C574,C577-C579|FallopianTube|911|Mesonephroma|9110/3|Mesonephroma
C571-C574,C577-C579|FallopianTube|959|Lymphoma|9590/3|Lymphoma
C571-C574,C577-C579|FallopianTube|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C571-C574,C577-C579|FallopianTube|959|Lymphoma|9596/3|CompositeLymphoma
C571-C574,C577-C579|FallopianTube|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C571-C574,C577-C579|FallopianTube|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C571-C574,C577-C579|FallopianTube|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C571-C574,C577-C579|FallopianTube|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C571-C574,C577-C579|FallopianTube|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C571-C574,C577-C579|FallopianTube|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C571-C574,C577-C579|FallopianTube|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C571-C574,C577-C579|FallopianTube|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C571-C574,C577-C579|FallopianTube|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C571-C574,C577-C579|FallopianTube|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C571-C574,C577-C579|FallopianTube|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C571-C574,C577-C579|FallopianTube|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C571-C574,C577-C579|FallopianTube|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C571-C574,C577-C579|FallopianTube|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C571-C574,C577-C579|FallopianTube|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C571-C574,C577-C579|FallopianTube|967|BCellLymphomas|9673/3|MantleCellLymphoma
C571-C574,C577-C579|FallopianTube|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C571-C574,C577-C579|FallopianTube|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C571-C574,C577-C579|FallopianTube|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C571-C574,C577-C579|FallopianTube|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C571-C574,C577-C579|FallopianTube|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C571-C574,C577-C579|FallopianTube|969|FollicularAdenoma|9690/3|LymphomaFollicular
C571-C574,C577-C579|FallopianTube|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C571-C574,C577-C579|FallopianTube|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C571-C574,C577-C579|FallopianTube|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C571-C574,C577-C579|FallopianTube|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C571-C574,C577-C579|FallopianTube|970|TCellLymphoma|9701/3|SezarySyndrome
C571-C574,C577-C579|FallopianTube|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C571-C574,C577-C579|FallopianTube|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C571-C574,C577-C579|FallopianTube|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C571-C574,C577-C579|FallopianTube|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C571-C574,C577-C579|FallopianTube|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C571-C574,C577-C579|FallopianTube|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C571-C574,C577-C579|FallopianTube|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C571-C574,C577-C579|FallopianTube|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C571-C574,C577-C579|FallopianTube|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C571-C574,C577-C579|FallopianTube|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C571-C574,C577-C579|FallopianTube|973|Plasmacytoma|9731/3|Plasmacytoma
C571-C574,C577-C579|FallopianTube|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C571-C574,C577-C579|FallopianTube|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C571-C574,C577-C579|FallopianTube|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C571-C574,C577-C579|FallopianTube|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C571-C574,C577-C579|FallopianTube|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C571-C574,C577-C579|FallopianTube|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C571-C574,C577-C579|FallopianTube|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C571-C574,C577-C579|FallopianTube|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C571-C574,C577-C579|FallopianTube|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C571-C574,C577-C579|FallopianTube|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C571-C574,C577-C579|FallopianTube|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C571-C574,C577-C579|FallopianTube|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C571-C574,C577-C579|FallopianTube|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C571-C574,C577-C579|FallopianTube|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C571-C574,C577-C579|FallopianTube|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C571-C574,C577-C579|FallopianTube|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9812/3|null
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9813/3|null
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9814/3|null
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9817/3|null
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9818/3|null
C571-C574,C577-C579|FallopianTube|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C571-C574,C577-C579|FallopianTube|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C571-C574,C577-C579|FallopianTube|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C571-C574,C577-C579|FallopianTube|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C571-C574,C577-C579|FallopianTube|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C571-C574,C577-C579|FallopianTube|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C571-C574,C577-C579|FallopianTube|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C571-C574,C577-C579|FallopianTube|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C589|PlacentaPart|910|Choriocarcinoma|9100/3|Choriocarcinoma
C589|PlacentaPart|910|Choriocarcinoma|9101/3|Choriocarcinoma
C589|PlacentaPart|910|Choriocarcinoma|9104/3|PlacentalSiteGTT
C589|PlacentaPart|910|Choriocarcinoma|9105/3|EpithelioidTrophoblasticTumor
C589|PlacentaPart|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C589|PlacentaPart|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C600-C602,C608-C609|Penis|801|Carcinoma|8010/2|InSituCancer
C600-C602,C608-C609|Penis|801|Carcinoma|8010/3|CarcinomaNOSDNE
C600-C602,C608-C609|Penis|801|Carcinoma|8011/3|MalignantEpithelioma
C600-C602,C608-C609|Penis|801|Carcinoma|8012/3|LargeCellCarcinoma
C600-C602,C608-C609|Penis|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C600-C602,C608-C609|Penis|801|Carcinoma|8014/3|LargeCellCarcinoma
C600-C602,C608-C609|Penis|801|Carcinoma|8015/3|GlassyCellCarcinoma
C600-C602,C608-C609|Penis|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C600-C602,C608-C609|Penis|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C600-C602,C608-C609|Penis|802|Carcinoma|8022/3|PleomorphicCarcinoma
C600-C602,C608-C609|Penis|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C600-C602,C608-C609|Penis|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C600-C602,C608-C609|Penis|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C600-C602,C608-C609|Penis|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C600-C602,C608-C609|Penis|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C600-C602,C608-C609|Penis|805|PapillaryCarcinoma|8054/3|VerrucousCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8071/2|KeratinizingSquamousCellCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C600-C602,C608-C609|Penis|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C600-C602,C608-C609|Penis|808|LymphoepithelialCarcinoma|8080/2|PenileCarcinomaInSitu
C600-C602,C608-C609|Penis|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C600-C602,C608-C609|Penis|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C600-C602,C608-C609|Penis|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C600-C602,C608-C609|Penis|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C600-C602,C608-C609|Penis|809|BasalCellCarcinoma|8090/3|BasalCellCarcinoma
C600-C602,C608-C609|Penis|809|BasalCellCarcinoma|8091/3|SuperficialBasalCellCarcinoma
C600-C602,C608-C609|Penis|809|BasalCellCarcinoma|8092/3|SkinInfiltratingBasalCellCarcinoma
C600-C602,C608-C609|Penis|809|BasalCellCarcinoma|8093/3|FibroepitheliomaOfPinkus
C600-C602,C608-C609|Penis|809|BasalCellCarcinoma|8094/3|SkinBasosquamousCellCarcinoma
C600-C602,C608-C609|Penis|809|BasalCellCarcinoma|8095/3|SkinMetatypicalCarcinoma
C600-C602,C608-C609|Penis|809|BasalCellCarcinoma|8097/3|SkinNodularBasalCellCarcinoma
C600-C602,C608-C609|Penis|809|BasalCellCarcinoma|8098/3|SkinAdenoidBasalCellCarcinoma
C600-C602,C608-C609|Penis|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C600-C602,C608-C609|Penis|811|PilomatricalCarcinoma|8110/3|PilomatricalCarcinoma
C600-C602,C608-C609|Penis|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C600-C602,C608-C609|Penis|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C600-C602,C608-C609|Penis|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C600-C602,C608-C609|Penis|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C600-C602,C608-C609|Penis|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C600-C602,C608-C609|Penis|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8140/3|Adenocarcinoma
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C600-C602,C608-C609|Penis|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C600-C602,C608-C609|Penis|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C600-C602,C608-C609|Penis|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C600-C602,C608-C609|Penis|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C600-C602,C608-C609|Penis|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C600-C602,C608-C609|Penis|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C600-C602,C608-C609|Penis|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C600-C602,C608-C609|Penis|839|AdnexalCarcinoma|8390/3|AdnexalCarcinoma
C600-C602,C608-C609|Penis|840|SweatGlandAdenocarcinoma|8400/3|SweatGlandAdenocarcinoma
C600-C602,C608-C609|Penis|840|SweatGlandAdenocarcinoma|8401/3|ApocrineAdenocarcinoma
C600-C602,C608-C609|Penis|841|EccrineAdenocarcinoma|8410/3|SebaceousAdenocarcinoma
C600-C602,C608-C609|Penis|841|EccrineAdenocarcinoma|8413/3|EccrineAdenocarcinoma
C600-C602,C608-C609|Penis|854|PagetDiseaseExtramammary|8542/3|PagetDiseaseExtramammary
C600-C602,C608-C609|Penis|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C600-C602,C608-C609|Penis|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C600-C602,C608-C609|Penis|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C600-C602,C608-C609|Penis|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C600-C602,C608-C609|Penis|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C600-C602,C608-C609|Penis|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C600-C602,C608-C609|Penis|872|Melanoma|8720/2|Stage0SkinMelanoma
C600-C602,C608-C609|Penis|872|Melanoma|8720/3|Melanoma
C600-C602,C608-C609|Penis|872|Melanoma|8721/3|NodularMelanoma
C600-C602,C608-C609|Penis|872|Melanoma|8722/3|BalloonCellMelanoma
C600-C602,C608-C609|Penis|872|Melanoma|8723/3|RegressingMelanoma
C600-C602,C608-C609|Penis|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C600-C602,C608-C609|Penis|874|Nevus|8740/3|MelanomaInJunctionalNevus
C600-C602,C608-C609|Penis|874|Nevus|8741/2|PrecancerousMelanosis
C600-C602,C608-C609|Penis|874|Nevus|8741/3|Melanoma
C600-C602,C608-C609|Penis|874|Nevus|8742/2|LentigoMaligna
C600-C602,C608-C609|Penis|874|Nevus|8742/3|LentigoMalignaMelanoma
C600-C602,C608-C609|Penis|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C600-C602,C608-C609|Penis|874|Nevus|8745/3|DesmoplasticMelanoma
C600-C602,C608-C609|Penis|874|Nevus|8746/3|MucosalLentiginousMelanoma
C600-C602,C608-C609|Penis|876|Nevus|8761/3|GiantCongenitalNevus
C600-C602,C608-C609|Penis|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C600-C602,C608-C609|Penis|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C600-C602,C608-C609|Penis|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C600-C602,C608-C609|Penis|878|MelanomaArisingFromBlueNevus|8780/3|MelanomaArisingFromBlueNevus
C600-C602,C608-C609|Penis|880|Sarcoma|8800/3|Sarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8801/3|SpindleCellSarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8802/3|GiantCellSarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8803/3|SmallCellSarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8804/3|SarcomaEpithelioid
C600-C602,C608-C609|Penis|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C600-C602,C608-C609|Penis|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C600-C602,C608-C609|Penis|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C600-C602,C608-C609|Penis|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C600-C602,C608-C609|Penis|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C600-C602,C608-C609|Penis|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C600-C602,C608-C609|Penis|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C600-C602,C608-C609|Penis|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8850/3|Liposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C600-C602,C608-C609|Penis|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8855/3|Liposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C600-C602,C608-C609|Penis|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C600-C602,C608-C609|Penis|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C600-C602,C608-C609|Penis|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C600-C602,C608-C609|Penis|889|MyomatousNeoplasm|8895/3|Myosarcoma
C600-C602,C608-C609|Penis|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C600-C602,C608-C609|Penis|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C600-C602,C608-C609|Penis|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C600-C602,C608-C609|Penis|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C600-C602,C608-C609|Penis|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C600-C602,C608-C609|Penis|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C600-C602,C608-C609|Penis|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C600-C602,C608-C609|Penis|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C600-C602,C608-C609|Penis|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C600-C602,C608-C609|Penis|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C600-C602,C608-C609|Penis|898|Carcinosarcoma|8980/3|Carcinosarcoma
C600-C602,C608-C609|Penis|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C600-C602,C608-C609|Penis|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C600-C602,C608-C609|Penis|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C600-C602,C608-C609|Penis|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C600-C602,C608-C609|Penis|914|KaposiSarcoma|9140/3|KaposiSarcoma
C600-C602,C608-C609|Penis|959|Lymphoma|9597/3|CrostisDisease
C600-C602,C608-C609|Penis|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C600-C602,C608-C609|Penis|970|TCellLymphoma|9700/3|MycosisFungoides
C600-C602,C608-C609|Penis|970|TCellLymphoma|9701/3|SezarySyndrome
C600-C602,C608-C609|Penis|970|TCellLymphoma|9708/3|TCellLymphoma
C600-C602,C608-C609|Penis|970|TCellLymphoma|9709/3|CutaneousTCellNonHodgkinLymphoma
C600-C602,C608-C609|Penis|971|AdultNonHodgkinLymphoma|9718/3|CALCL
C600-C602,C608-C609|Penis|972|LymphoblasticLymphoma|9725/3|HydroaVacciniformeLikeLymphoma
C600-C602,C608-C609|Penis|972|LymphoblasticLymphoma|9726/3|TCellLymphoma
C600-C602,C608-C609|Penis|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C619|Prostate|801|Carcinoma|8010/2|InSituCancer
C619|Prostate|801|Carcinoma|8010/3|CarcinomaNOSDNE
C619|Prostate|801|Carcinoma|8011/3|MalignantEpithelioma
C619|Prostate|801|Carcinoma|8012/3|LargeCellCarcinoma
C619|Prostate|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C619|Prostate|801|Carcinoma|8014/3|LargeCellCarcinoma
C619|Prostate|801|Carcinoma|8015/3|GlassyCellCarcinoma
C619|Prostate|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C619|Prostate|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C619|Prostate|802|Carcinoma|8022/3|PleomorphicCarcinoma
C619|Prostate|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C619|Prostate|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C619|Prostate|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C619|Prostate|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C619|Prostate|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C619|Prostate|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C619|Prostate|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C619|Prostate|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C619|Prostate|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C619|Prostate|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C619|Prostate|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C619|Prostate|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C619|Prostate|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C619|Prostate|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C619|Prostate|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C619|Prostate|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C619|Prostate|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C619|Prostate|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C619|Prostate|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C619|Prostate|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C619|Prostate|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C619|Prostate|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C619|Prostate|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C619|Prostate|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C619|Prostate|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C619|Prostate|814|Adenocarcinoma|8140/1|MalignantProstateNeoplasm
C619|Prostate|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C619|Prostate|814|Adenocarcinoma|8140/3|Adenocarcinoma
C619|Prostate|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C619|Prostate|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C619|Prostate|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C619|Prostate|814|Adenocarcinoma|8148/2|IntraepithelialNeoplasia
C619|Prostate|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C619|Prostate|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C619|Prostate|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C619|Prostate|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C619|Prostate|825|BronchioloalveolarAdenocarcinoma|8251/3|BronchioloalveolarAdenocarcinoma
C619|Prostate|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C619|Prostate|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C619|Prostate|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C619|Prostate|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C619|Prostate|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C619|Prostate|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C619|Prostate|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C619|Prostate|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C619|Prostate|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C619|Prostate|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C619|Prostate|850|DuctalCarcinoma|8500/2|DuctalBreastCarcinomaInSitu
C619|Prostate|850|DuctalCarcinoma|8500/3|InvasiveBreastCarcinoma
C619|Prostate|850|DuctalCarcinoma|8503/2|IntraductalPapillaryBreastCarcinoma
C619|Prostate|850|DuctalCarcinoma|8503/3|IntraductalPapillaryBreastCarcinoma
C619|Prostate|850|DuctalCarcinoma|8504/2|IntracysticPapillaryBreastCarcinoma
C619|Prostate|850|DuctalCarcinoma|8504/3|IntracysticPapillaryBreastCarcinoma
C619|Prostate|850|DuctalCarcinoma|8507/2|MicropapillaryCarcinoma
C619|Prostate|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C619|Prostate|851|MedullaryCarcinoma|8514/3|DesmoplasticNodularMedulloblastoma
C619|Prostate|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C619|Prostate|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C619|Prostate|855|AcinarCellCarcinoma|8552/3|ProstateAcinarAdenocarcinoma
C619|Prostate|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C619|Prostate|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C619|Prostate|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C619|Prostate|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C619|Prostate|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C619|Prostate|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C619|Prostate|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C619|Prostate|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C619|Prostate|880|Sarcoma|8800/3|Sarcoma
C619|Prostate|880|Sarcoma|8801/3|SpindleCellSarcoma
C619|Prostate|880|Sarcoma|8802/3|GiantCellSarcoma
C619|Prostate|880|Sarcoma|8803/3|SmallCellSarcoma
C619|Prostate|880|Sarcoma|8804/3|SarcomaEpithelioid
C619|Prostate|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C619|Prostate|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C619|Prostate|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C619|Prostate|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C619|Prostate|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C619|Prostate|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C619|Prostate|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C619|Prostate|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C619|Prostate|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C619|Prostate|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C619|Prostate|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C619|Prostate|889|MyomatousNeoplasm|8895/3|Myosarcoma
C619|Prostate|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C619|Prostate|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C619|Prostate|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C619|Prostate|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C619|Prostate|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C619|Prostate|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C619|Prostate|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C619|Prostate|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C619|Prostate|898|Carcinosarcoma|8980/3|Carcinosarcoma
C619|Prostate|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C619|Prostate|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C619|Prostate|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C619|Prostate|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C619|Prostate|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C619|Prostate|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C619|Prostate|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C619|Prostate|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C619|Prostate|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C619|Prostate|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C619|Prostate|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C619|Prostate|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C619|Prostate|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C619|Prostate|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C619|Prostate|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C619|Prostate|981|PrecursorLymphoidNeoplasm|9812/3|null
C619|Prostate|981|PrecursorLymphoidNeoplasm|9813/3|null
C619|Prostate|981|PrecursorLymphoidNeoplasm|9814/3|null
C619|Prostate|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C619|Prostate|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C619|Prostate|981|PrecursorLymphoidNeoplasm|9817/3|null
C619|Prostate|981|PrecursorLymphoidNeoplasm|9818/3|null
C619|Prostate|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C619|Prostate|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C619|Prostate|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C619|Prostate|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C619|Prostate|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C619|Prostate|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C619|Prostate|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C619|Prostate|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C620-C621,C629|Testis|801|Carcinoma|8010/2|InSituCancer
C620-C621,C629|Testis|801|Carcinoma|8010/3|CarcinomaNOSDNE
C620-C621,C629|Testis|801|Carcinoma|8011/3|MalignantEpithelioma
C620-C621,C629|Testis|801|Carcinoma|8012/3|LargeCellCarcinoma
C620-C621,C629|Testis|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C620-C621,C629|Testis|801|Carcinoma|8014/3|LargeCellCarcinoma
C620-C621,C629|Testis|801|Carcinoma|8015/3|GlassyCellCarcinoma
C620-C621,C629|Testis|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C620-C621,C629|Testis|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C620-C621,C629|Testis|802|Carcinoma|8022/3|PleomorphicCarcinoma
C620-C621,C629|Testis|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C620-C621,C629|Testis|814|Adenocarcinoma|8140/3|Adenocarcinoma
C620-C621,C629|Testis|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C620-C621,C629|Testis|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C620-C621,C629|Testis|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C620-C621,C629|Testis|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C620-C621,C629|Testis|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C620-C621,C629|Testis|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C620-C621,C629|Testis|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C620-C621,C629|Testis|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C620-C621,C629|Testis|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C620-C621,C629|Testis|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C620-C621,C629|Testis|863|GonadalNeoplasm|8630/3|MalignantSertoliCellTumor
C620-C621,C629|Testis|863|GonadalNeoplasm|8631/3|SertoliLeydigCellTumor
C620-C621,C629|Testis|863|GonadalNeoplasm|8634/3|SertoliLeydigCellTumor
C620-C621,C629|Testis|864|SertoliCellCarcinoma|8640/3|SertoliCellCarcinoma
C620-C621,C629|Testis|865|MalignantLeydigCellTumor|8650/3|MalignantLeydigCellTumor
C620-C621,C629|Testis|880|Sarcoma|8800/3|Sarcoma
C620-C621,C629|Testis|880|Sarcoma|8801/3|SpindleCellSarcoma
C620-C621,C629|Testis|880|Sarcoma|8802/3|GiantCellSarcoma
C620-C621,C629|Testis|880|Sarcoma|8803/3|SmallCellSarcoma
C620-C621,C629|Testis|880|Sarcoma|8804/3|SarcomaEpithelioid
C620-C621,C629|Testis|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C620-C621,C629|Testis|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C620-C621,C629|Testis|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C620-C621,C629|Testis|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C620-C621,C629|Testis|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C620-C621,C629|Testis|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C620-C621,C629|Testis|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C620-C621,C629|Testis|906|GermCellTumor|9060/3|Dysgerminoma
C620-C621,C629|Testis|906|GermCellTumor|9061/3|Seminoma
C620-C621,C629|Testis|906|GermCellTumor|9062/3|AtypicalSeminoma
C620-C621,C629|Testis|906|GermCellTumor|9063/3|TesticularSpermatocyticSeminoma
C620-C621,C629|Testis|906|GermCellTumor|9064/2|IntratubularGermCellNeoplasia
C620-C621,C629|Testis|906|GermCellTumor|9064/3|Germinoma
C620-C621,C629|Testis|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C620-C621,C629|Testis|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C620-C621,C629|Testis|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C620-C621,C629|Testis|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C620-C621,C629|Testis|908|Teratoma|9080/3|ImmatureTeratoma
C620-C621,C629|Testis|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C620-C621,C629|Testis|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C620-C621,C629|Testis|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C620-C621,C629|Testis|908|Teratoma|9084/3|Teratoma
C620-C621,C629|Testis|908|Teratoma|9085/3|MixedGermCellTumor
C620-C621,C629|Testis|910|Choriocarcinoma|9100/3|Choriocarcinoma
C620-C621,C629|Testis|910|Choriocarcinoma|9101/3|Choriocarcinoma
C620-C621,C629|Testis|910|Choriocarcinoma|9102/3|MalignantTrophoblasticTeratoma
C620-C621,C629|Testis|910|Choriocarcinoma|9105/3|EpithelioidTrophoblasticTumor
C620-C621,C629|Testis|959|Lymphoma|9590/3|Lymphoma
C620-C621,C629|Testis|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C620-C621,C629|Testis|959|Lymphoma|9596/3|CompositeLymphoma
C620-C621,C629|Testis|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C620-C621,C629|Testis|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C620-C621,C629|Testis|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C620-C621,C629|Testis|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C620-C621,C629|Testis|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C620-C621,C629|Testis|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C620-C621,C629|Testis|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C620-C621,C629|Testis|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C620-C621,C629|Testis|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C620-C621,C629|Testis|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C620-C621,C629|Testis|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C620-C621,C629|Testis|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C620-C621,C629|Testis|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C620-C621,C629|Testis|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C620-C621,C629|Testis|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C620-C621,C629|Testis|967|BCellLymphomas|9673/3|MantleCellLymphoma
C620-C621,C629|Testis|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C620-C621,C629|Testis|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C620-C621,C629|Testis|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C620-C621,C629|Testis|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C620-C621,C629|Testis|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C620-C621,C629|Testis|969|FollicularAdenoma|9690/3|LymphomaFollicular
C620-C621,C629|Testis|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C620-C621,C629|Testis|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C620-C621,C629|Testis|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C620-C621,C629|Testis|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C620-C621,C629|Testis|970|TCellLymphoma|9701/3|SezarySyndrome
C620-C621,C629|Testis|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C620-C621,C629|Testis|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C620-C621,C629|Testis|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C620-C621,C629|Testis|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C620-C621,C629|Testis|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C620-C621,C629|Testis|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C620-C621,C629|Testis|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C620-C621,C629|Testis|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C620-C621,C629|Testis|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C620-C621,C629|Testis|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C620-C621,C629|Testis|973|Plasmacytoma|9731/3|Plasmacytoma
C620-C621,C629|Testis|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C620-C621,C629|Testis|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C620-C621,C629|Testis|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C620-C621,C629|Testis|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C620-C621,C629|Testis|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C620-C621,C629|Testis|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C620-C621,C629|Testis|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C620-C621,C629|Testis|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C620-C621,C629|Testis|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C620-C621,C629|Testis|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C620-C621,C629|Testis|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C620-C621,C629|Testis|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C620-C621,C629|Testis|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C620-C621,C629|Testis|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C620-C621,C629|Testis|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C620-C621,C629|Testis|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9812/3|null
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9813/3|null
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9814/3|null
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9817/3|null
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9818/3|null
C620-C621,C629|Testis|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C620-C621,C629|Testis|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C620-C621,C629|Testis|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C620-C621,C629|Testis|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C620-C621,C629|Testis|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C620-C621,C629|Testis|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C620-C621,C629|Testis|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C620-C621,C629|Testis|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C630, C631, C637-C639|SpermaticCord|801|Carcinoma|8010/2|InSituCancer
C630, C631, C637-C639|SpermaticCord|801|Carcinoma|8010/3|CarcinomaNOSDNE
C630, C631, C637-C639|SpermaticCord|801|Carcinoma|8011/3|MalignantEpithelioma
C630, C631, C637-C639|SpermaticCord|801|Carcinoma|8012/3|LargeCellCarcinoma
C630, C631, C637-C639|SpermaticCord|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C630, C631, C637-C639|SpermaticCord|801|Carcinoma|8014/3|LargeCellCarcinoma
C630, C631, C637-C639|SpermaticCord|801|Carcinoma|8015/3|GlassyCellCarcinoma
C630, C631, C637-C639|SpermaticCord|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C630, C631, C637-C639|SpermaticCord|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C630, C631, C637-C639|SpermaticCord|802|Carcinoma|8022/3|PleomorphicCarcinoma
C630, C631, C637-C639|SpermaticCord|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C630, C631, C637-C639|SpermaticCord|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C630, C631, C637-C639|SpermaticCord|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C630, C631, C637-C639|SpermaticCord|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C630, C631, C637-C639|SpermaticCord|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C630, C631, C637-C639|SpermaticCord|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C630, C631, C637-C639|SpermaticCord|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C630, C631, C637-C639|SpermaticCord|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C630, C631, C637-C639|SpermaticCord|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C630, C631, C637-C639|SpermaticCord|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C630, C631, C637-C639|SpermaticCord|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C630, C631, C637-C639|SpermaticCord|814|Adenocarcinoma|8140/3|Adenocarcinoma
C630, C631, C637-C639|SpermaticCord|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C630, C631, C637-C639|SpermaticCord|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C630, C631, C637-C639|SpermaticCord|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C630, C631, C637-C639|SpermaticCord|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C630, C631, C637-C639|SpermaticCord|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C630, C631, C637-C639|SpermaticCord|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C630, C631, C637-C639|SpermaticCord|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C630, C631, C637-C639|SpermaticCord|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C630, C631, C637-C639|SpermaticCord|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C630, C631, C637-C639|SpermaticCord|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C630, C631, C637-C639|SpermaticCord|840|SweatGlandAdenocarcinoma|8401/3|ApocrineAdenocarcinoma
C630, C631, C637-C639|SpermaticCord|854|PagetDiseaseExtramammary|8542/3|PagetDiseaseExtramammary
C630, C631, C637-C639|SpermaticCord|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C630, C631, C637-C639|SpermaticCord|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C630, C631, C637-C639|SpermaticCord|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C630, C631, C637-C639|SpermaticCord|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C630, C631, C637-C639|SpermaticCord|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C630, C631, C637-C639|SpermaticCord|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C630, C631, C637-C639|SpermaticCord|880|Sarcoma|8800/3|Sarcoma
C630, C631, C637-C639|SpermaticCord|880|Sarcoma|8801/3|SpindleCellSarcoma
C630, C631, C637-C639|SpermaticCord|880|Sarcoma|8802/3|GiantCellSarcoma
C630, C631, C637-C639|SpermaticCord|880|Sarcoma|8803/3|SmallCellSarcoma
C630, C631, C637-C639|SpermaticCord|880|Sarcoma|8804/3|SarcomaEpithelioid
C630, C631, C637-C639|SpermaticCord|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C630, C631, C637-C639|SpermaticCord|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C630, C631, C637-C639|SpermaticCord|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C630, C631, C637-C639|SpermaticCord|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C630, C631, C637-C639|SpermaticCord|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C630, C631, C637-C639|SpermaticCord|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C630, C631, C637-C639|SpermaticCord|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C630, C631, C637-C639|SpermaticCord|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C630, C631, C637-C639|SpermaticCord|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C630, C631, C637-C639|SpermaticCord|885|Liposarcoma|8850/3|Liposarcoma
C630, C631, C637-C639|SpermaticCord|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C630, C631, C637-C639|SpermaticCord|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C630, C631, C637-C639|SpermaticCord|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C630, C631, C637-C639|SpermaticCord|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C630, C631, C637-C639|SpermaticCord|885|Liposarcoma|8855/3|Liposarcoma
C630, C631, C637-C639|SpermaticCord|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C630, C631, C637-C639|SpermaticCord|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C630, C631, C637-C639|SpermaticCord|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C630, C631, C637-C639|SpermaticCord|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C630, C631, C637-C639|SpermaticCord|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C630, C631, C637-C639|SpermaticCord|889|MyomatousNeoplasm|8895/3|Myosarcoma
C630, C631, C637-C639|SpermaticCord|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C630, C631, C637-C639|SpermaticCord|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C630, C631, C637-C639|SpermaticCord|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C630, C631, C637-C639|SpermaticCord|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C630, C631, C637-C639|SpermaticCord|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C630, C631, C637-C639|SpermaticCord|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C630, C631, C637-C639|SpermaticCord|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C630, C631, C637-C639|SpermaticCord|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C630, C631, C637-C639|SpermaticCord|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C630, C631, C637-C639|SpermaticCord|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C630, C631, C637-C639|SpermaticCord|898|Carcinosarcoma|8980/3|Carcinosarcoma
C630, C631, C637-C639|SpermaticCord|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C630, C631, C637-C639|SpermaticCord|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C630, C631, C637-C639|SpermaticCord|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C630, C631, C637-C639|SpermaticCord|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C630, C631, C637-C639|SpermaticCord|914|KaposiSarcoma|9140/3|KaposiSarcoma
C630, C631, C637-C639|SpermaticCord|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C630, C631, C637-C639|SpermaticCord|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C632|Scrotum|801|Carcinoma|8010/2|InSituCancer
C632|Scrotum|801|Carcinoma|8010/3|CarcinomaNOSDNE
C632|Scrotum|801|Carcinoma|8011/3|MalignantEpithelioma
C632|Scrotum|801|Carcinoma|8012/3|LargeCellCarcinoma
C632|Scrotum|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C632|Scrotum|801|Carcinoma|8014/3|LargeCellCarcinoma
C632|Scrotum|801|Carcinoma|8015/3|GlassyCellCarcinoma
C632|Scrotum|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C632|Scrotum|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C632|Scrotum|802|Carcinoma|8022/3|PleomorphicCarcinoma
C632|Scrotum|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C632|Scrotum|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C632|Scrotum|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C632|Scrotum|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C632|Scrotum|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C632|Scrotum|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C632|Scrotum|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C632|Scrotum|808|LymphoepithelialCarcinoma|8080/2|PenileCarcinomaInSitu
C632|Scrotum|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C632|Scrotum|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C632|Scrotum|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C632|Scrotum|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C632|Scrotum|809|BasalCellCarcinoma|8090/3|BasalCellCarcinoma
C632|Scrotum|809|BasalCellCarcinoma|8091/3|SuperficialBasalCellCarcinoma
C632|Scrotum|809|BasalCellCarcinoma|8092/3|SkinInfiltratingBasalCellCarcinoma
C632|Scrotum|809|BasalCellCarcinoma|8093/3|FibroepitheliomaOfPinkus
C632|Scrotum|809|BasalCellCarcinoma|8094/3|SkinBasosquamousCellCarcinoma
C632|Scrotum|809|BasalCellCarcinoma|8095/3|SkinMetatypicalCarcinoma
C632|Scrotum|809|BasalCellCarcinoma|8097/3|SkinNodularBasalCellCarcinoma
C632|Scrotum|809|BasalCellCarcinoma|8098/3|SkinAdenoidBasalCellCarcinoma
C632|Scrotum|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C632|Scrotum|811|PilomatricalCarcinoma|8110/3|PilomatricalCarcinoma
C632|Scrotum|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C632|Scrotum|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C632|Scrotum|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C632|Scrotum|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C632|Scrotum|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C632|Scrotum|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C632|Scrotum|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C632|Scrotum|814|Adenocarcinoma|8140/3|Adenocarcinoma
C632|Scrotum|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C632|Scrotum|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C632|Scrotum|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C632|Scrotum|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C632|Scrotum|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C632|Scrotum|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C632|Scrotum|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C632|Scrotum|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C632|Scrotum|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C632|Scrotum|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C632|Scrotum|839|AdnexalCarcinoma|8390/3|AdnexalCarcinoma
C632|Scrotum|840|SweatGlandAdenocarcinoma|8400/3|SweatGlandAdenocarcinoma
C632|Scrotum|840|SweatGlandAdenocarcinoma|8401/3|ApocrineAdenocarcinoma
C632|Scrotum|841|EccrineAdenocarcinoma|8410/3|SebaceousAdenocarcinoma
C632|Scrotum|841|EccrineAdenocarcinoma|8413/3|EccrineAdenocarcinoma
C632|Scrotum|854|PagetDiseaseExtramammary|8542/3|PagetDiseaseExtramammary
C632|Scrotum|857|AdenocarcinomaWithMetaplasia|8570/3|AdenocarcinomaWithSquamousMetaplasia
C632|Scrotum|857|AdenocarcinomaWithMetaplasia|8571/3|AdenocarcinomaWithOsseousMetaplasia
C632|Scrotum|857|AdenocarcinomaWithMetaplasia|8572/3|AdenocarcinomaSpindleCell
C632|Scrotum|857|AdenocarcinomaWithMetaplasia|8573/3|AdenocarcinomaWithApocrineMetaplasia
C632|Scrotum|857|AdenocarcinomaWithMetaplasia|8574/3|NeuroendocrineNeoplasm
C632|Scrotum|857|AdenocarcinomaWithMetaplasia|8575/3|MetaplasticCarcinoma
C632|Scrotum|872|Melanoma|8720/2|Stage0SkinMelanoma
C632|Scrotum|872|Melanoma|8720/3|Melanoma
C632|Scrotum|872|Melanoma|8721/3|NodularMelanoma
C632|Scrotum|872|Melanoma|8722/3|BalloonCellMelanoma
C632|Scrotum|872|Melanoma|8723/3|RegressingMelanoma
C632|Scrotum|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C632|Scrotum|874|Nevus|8740/3|MelanomaInJunctionalNevus
C632|Scrotum|874|Nevus|8741/2|PrecancerousMelanosis
C632|Scrotum|874|Nevus|8741/3|Melanoma
C632|Scrotum|874|Nevus|8742/2|LentigoMaligna
C632|Scrotum|874|Nevus|8742/3|LentigoMalignaMelanoma
C632|Scrotum|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C632|Scrotum|874|Nevus|8745/3|DesmoplasticMelanoma
C632|Scrotum|874|Nevus|8746/3|MucosalLentiginousMelanoma
C632|Scrotum|876|Nevus|8761/3|GiantCongenitalNevus
C632|Scrotum|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C632|Scrotum|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C632|Scrotum|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C632|Scrotum|878|MelanomaArisingFromBlueNevus|8780/3|MelanomaArisingFromBlueNevus
C632|Scrotum|880|Sarcoma|8800/3|Sarcoma
C632|Scrotum|880|Sarcoma|8801/3|SpindleCellSarcoma
C632|Scrotum|880|Sarcoma|8802/3|GiantCellSarcoma
C632|Scrotum|880|Sarcoma|8803/3|SmallCellSarcoma
C632|Scrotum|880|Sarcoma|8804/3|SarcomaEpithelioid
C632|Scrotum|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C632|Scrotum|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C632|Scrotum|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C632|Scrotum|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C632|Scrotum|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C632|Scrotum|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C632|Scrotum|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C632|Scrotum|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C632|Scrotum|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C632|Scrotum|885|Liposarcoma|8850/3|Liposarcoma
C632|Scrotum|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C632|Scrotum|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C632|Scrotum|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C632|Scrotum|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C632|Scrotum|885|Liposarcoma|8855/3|Liposarcoma
C632|Scrotum|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C632|Scrotum|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C632|Scrotum|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C632|Scrotum|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C632|Scrotum|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C632|Scrotum|889|MyomatousNeoplasm|8895/3|Myosarcoma
C632|Scrotum|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C632|Scrotum|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C632|Scrotum|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C632|Scrotum|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C632|Scrotum|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C632|Scrotum|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C632|Scrotum|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C632|Scrotum|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C632|Scrotum|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C632|Scrotum|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C632|Scrotum|898|Carcinosarcoma|8980/3|Carcinosarcoma
C632|Scrotum|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C632|Scrotum|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C632|Scrotum|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C632|Scrotum|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C632|Scrotum|914|KaposiSarcoma|9140/3|KaposiSarcoma
C632|Scrotum|959|Lymphoma|9597/3|CrostisDisease
C632|Scrotum|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C632|Scrotum|970|TCellLymphoma|9700/3|MycosisFungoides
C632|Scrotum|970|TCellLymphoma|9701/3|SezarySyndrome
C632|Scrotum|970|TCellLymphoma|9708/3|TCellLymphoma
C632|Scrotum|970|TCellLymphoma|9709/3|CutaneousTCellNonHodgkinLymphoma
C632|Scrotum|971|AdultNonHodgkinLymphoma|9718/3|CALCL
C632|Scrotum|972|LymphoblasticLymphoma|9725/3|HydroaVacciniformeLikeLymphoma
C632|Scrotum|972|LymphoblasticLymphoma|9726/3|TCellLymphoma
C632|Scrotum|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C649|Kidney|801|Carcinoma|8010/2|InSituCancer
C649|Kidney|801|Carcinoma|8010/3|CarcinomaNOSDNE
C649|Kidney|801|Carcinoma|8011/3|MalignantEpithelioma
C649|Kidney|801|Carcinoma|8012/3|LargeCellCarcinoma
C649|Kidney|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C649|Kidney|801|Carcinoma|8014/3|LargeCellCarcinoma
C649|Kidney|801|Carcinoma|8015/3|GlassyCellCarcinoma
C649|Kidney|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C649|Kidney|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C649|Kidney|802|Carcinoma|8022/3|PleomorphicCarcinoma
C649|Kidney|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C649|Kidney|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C649|Kidney|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C649|Kidney|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C649|Kidney|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C649|Kidney|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C649|Kidney|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C649|Kidney|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C649|Kidney|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C649|Kidney|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C649|Kidney|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C649|Kidney|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C649|Kidney|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C649|Kidney|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C649|Kidney|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C649|Kidney|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C649|Kidney|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C649|Kidney|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C649|Kidney|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C649|Kidney|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C649|Kidney|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C649|Kidney|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C649|Kidney|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C649|Kidney|813|PapillaryTransitionalCellCarcinoma|8130/3|PapillaryTransitionalCellCarcinoma
C649|Kidney|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C649|Kidney|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C649|Kidney|814|Adenocarcinoma|8140/3|Adenocarcinoma
C649|Kidney|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C649|Kidney|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C649|Kidney|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C649|Kidney|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C649|Kidney|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C649|Kidney|823|SolidCarcinoma|8230/2|InSituCancer
C649|Kidney|823|SolidCarcinoma|8230/3|SolidCarcinoma
C649|Kidney|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C649|Kidney|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C649|Kidney|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C649|Kidney|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C649|Kidney|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C649|Kidney|831|ClearCellAdenocarcinoma|8311/3|RenalCellCarcinoma
C649|Kidney|831|ClearCellAdenocarcinoma|8312/3|RenalCellCarcinoma
C649|Kidney|831|ClearCellAdenocarcinoma|8316/3|CystassociatedRenalCellCarcinoma
C649|Kidney|831|ClearCellAdenocarcinoma|8317/3|ChromophobeRenalCellCarcinoma
C649|Kidney|831|ClearCellAdenocarcinoma|8318/3|SarcomatoidRenalCellCarcinoma
C649|Kidney|831|ClearCellAdenocarcinoma|8319/3|CollectingDuctCarcinomaOfKidney
C649|Kidney|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C649|Kidney|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C649|Kidney|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C649|Kidney|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C649|Kidney|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C649|Kidney|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C649|Kidney|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C649|Kidney|880|Sarcoma|8800/3|Sarcoma
C649|Kidney|880|Sarcoma|8801/3|SpindleCellSarcoma
C649|Kidney|880|Sarcoma|8802/3|GiantCellSarcoma
C649|Kidney|880|Sarcoma|8803/3|SmallCellSarcoma
C649|Kidney|880|Sarcoma|8804/3|SarcomaEpithelioid
C649|Kidney|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C649|Kidney|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C649|Kidney|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C649|Kidney|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C649|Kidney|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C649|Kidney|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C649|Kidney|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C649|Kidney|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C649|Kidney|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C649|Kidney|885|Liposarcoma|8850/3|Liposarcoma
C649|Kidney|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C649|Kidney|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C649|Kidney|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C649|Kidney|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C649|Kidney|885|Liposarcoma|8855/3|Liposarcoma
C649|Kidney|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C649|Kidney|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C649|Kidney|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C649|Kidney|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C649|Kidney|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C649|Kidney|889|MyomatousNeoplasm|8895/3|Myosarcoma
C649|Kidney|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C649|Kidney|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C649|Kidney|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C649|Kidney|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C649|Kidney|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C649|Kidney|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C649|Kidney|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C649|Kidney|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C649|Kidney|895|MixedTumorMullerian|8959/3|MalignantCysticNephroma
C649|Kidney|896|Nephroblastoma|8960/3|Nephroblastoma
C649|Kidney|896|Nephroblastoma|8963/3|RhabdoidTumor
C649|Kidney|896|Nephroblastoma|8964/3|ClearCellSarcomaOfTheKidney
C649|Kidney|898|Carcinosarcoma|8980/3|Carcinosarcoma
C649|Kidney|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C649|Kidney|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C649|Kidney|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C649|Kidney|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C649|Kidney|950|Neuroblastoma|9500/3|Neuroblastoma
C649|Kidney|950|Neuroblastoma|9501/3|Medulloepithelioma
C649|Kidney|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C649|Kidney|950|Neuroblastoma|9503/3|Neuroepithelioma
C649|Kidney|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C649|Kidney|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C649|Kidney|959|Lymphoma|9590/3|Lymphoma
C649|Kidney|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C649|Kidney|959|Lymphoma|9596/3|CompositeLymphoma
C649|Kidney|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C649|Kidney|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C649|Kidney|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C649|Kidney|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C649|Kidney|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C649|Kidney|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C649|Kidney|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C649|Kidney|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C649|Kidney|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C649|Kidney|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C649|Kidney|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C649|Kidney|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C649|Kidney|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C649|Kidney|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C649|Kidney|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C649|Kidney|967|BCellLymphomas|9673/3|MantleCellLymphoma
C649|Kidney|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C649|Kidney|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C649|Kidney|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C649|Kidney|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C649|Kidney|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C649|Kidney|969|FollicularAdenoma|9690/3|LymphomaFollicular
C649|Kidney|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C649|Kidney|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C649|Kidney|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C649|Kidney|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C649|Kidney|970|TCellLymphoma|9701/3|SezarySyndrome
C649|Kidney|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C649|Kidney|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C649|Kidney|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C649|Kidney|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C649|Kidney|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C649|Kidney|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C649|Kidney|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C649|Kidney|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C649|Kidney|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C649|Kidney|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C649|Kidney|973|Plasmacytoma|9731/3|Plasmacytoma
C649|Kidney|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C649|Kidney|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C649|Kidney|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C649|Kidney|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C649|Kidney|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C649|Kidney|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C649|Kidney|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C649|Kidney|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C649|Kidney|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C649|Kidney|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C649|Kidney|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C649|Kidney|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C649|Kidney|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C649|Kidney|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C649|Kidney|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C649|Kidney|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C649|Kidney|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C649|Kidney|981|PrecursorLymphoidNeoplasm|9812/3|null
C649|Kidney|981|PrecursorLymphoidNeoplasm|9813/3|null
C649|Kidney|981|PrecursorLymphoidNeoplasm|9814/3|null
C649|Kidney|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C649|Kidney|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C649|Kidney|981|PrecursorLymphoidNeoplasm|9817/3|null
C649|Kidney|981|PrecursorLymphoidNeoplasm|9818/3|null
C649|Kidney|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C649|Kidney|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C649|Kidney|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C649|Kidney|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C649|Kidney|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C649|Kidney|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C649|Kidney|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C649|Kidney|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C659, C669|RenalPelvis|801|Carcinoma|8010/2|InSituCancer
C659, C669|RenalPelvis|801|Carcinoma|8010/3|CarcinomaNOSDNE
C659, C669|RenalPelvis|801|Carcinoma|8011/3|MalignantEpithelioma
C659, C669|RenalPelvis|801|Carcinoma|8012/3|LargeCellCarcinoma
C659, C669|RenalPelvis|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C659, C669|RenalPelvis|801|Carcinoma|8014/3|LargeCellCarcinoma
C659, C669|RenalPelvis|801|Carcinoma|8015/3|GlassyCellCarcinoma
C659, C669|RenalPelvis|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C659, C669|RenalPelvis|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C659, C669|RenalPelvis|802|Carcinoma|8022/3|PleomorphicCarcinoma
C659, C669|RenalPelvis|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C659, C669|RenalPelvis|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C659, C669|RenalPelvis|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C659, C669|RenalPelvis|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C659, C669|RenalPelvis|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C659, C669|RenalPelvis|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C659, C669|RenalPelvis|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C659, C669|RenalPelvis|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C659, C669|RenalPelvis|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C659, C669|RenalPelvis|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C659, C669|RenalPelvis|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C659, C669|RenalPelvis|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C659, C669|RenalPelvis|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C659, C669|RenalPelvis|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C659, C669|RenalPelvis|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C659, C669|RenalPelvis|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C659, C669|RenalPelvis|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C659, C669|RenalPelvis|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C659, C669|RenalPelvis|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C659, C669|RenalPelvis|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C659, C669|RenalPelvis|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C659, C669|RenalPelvis|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C659, C669|RenalPelvis|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C659, C669|RenalPelvis|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C659, C669|RenalPelvis|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C659, C669|RenalPelvis|814|Adenocarcinoma|8140/3|Adenocarcinoma
C659, C669|RenalPelvis|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C659, C669|RenalPelvis|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C659, C669|RenalPelvis|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C659, C669|RenalPelvis|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C659, C669|RenalPelvis|821|AdenocarcinomaInAdenomatousPolyp|8211/3|TubularAdenocarcinoma
C659, C669|RenalPelvis|823|SolidCarcinoma|8230/2|InSituCancer
C659, C669|RenalPelvis|823|SolidCarcinoma|8230/3|SolidCarcinoma
C659, C669|RenalPelvis|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C659, C669|RenalPelvis|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C659, C669|RenalPelvis|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C659, C669|RenalPelvis|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C659, C669|RenalPelvis|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C659, C669|RenalPelvis|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C659, C669|RenalPelvis|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C659, C669|RenalPelvis|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C659, C669|RenalPelvis|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C659, C669|RenalPelvis|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C659, C669|RenalPelvis|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C659, C669|RenalPelvis|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C659, C669|RenalPelvis|880|Sarcoma|8800/3|Sarcoma
C659, C669|RenalPelvis|880|Sarcoma|8801/3|SpindleCellSarcoma
C659, C669|RenalPelvis|880|Sarcoma|8802/3|GiantCellSarcoma
C659, C669|RenalPelvis|880|Sarcoma|8803/3|SmallCellSarcoma
C659, C669|RenalPelvis|880|Sarcoma|8804/3|SarcomaEpithelioid
C659, C669|RenalPelvis|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C659, C669|RenalPelvis|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C659, C669|RenalPelvis|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C659, C669|RenalPelvis|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C659, C669|RenalPelvis|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C659, C669|RenalPelvis|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C659, C669|RenalPelvis|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C659, C669|RenalPelvis|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C659, C669|RenalPelvis|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C659, C669|RenalPelvis|885|Liposarcoma|8850/3|Liposarcoma
C659, C669|RenalPelvis|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C659, C669|RenalPelvis|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C659, C669|RenalPelvis|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C659, C669|RenalPelvis|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C659, C669|RenalPelvis|885|Liposarcoma|8855/3|Liposarcoma
C659, C669|RenalPelvis|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C659, C669|RenalPelvis|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C659, C669|RenalPelvis|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C659, C669|RenalPelvis|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C659, C669|RenalPelvis|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C659, C669|RenalPelvis|889|MyomatousNeoplasm|8895/3|Myosarcoma
C659, C669|RenalPelvis|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C659, C669|RenalPelvis|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C659, C669|RenalPelvis|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C659, C669|RenalPelvis|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C659, C669|RenalPelvis|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C659, C669|RenalPelvis|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C659, C669|RenalPelvis|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C659, C669|RenalPelvis|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C659, C669|RenalPelvis|895|MixedTumorMullerian|8959/3|MalignantCysticNephroma
C659, C669|RenalPelvis|896|Nephroblastoma|8964/3|ClearCellSarcomaOfTheKidney
C659, C669|RenalPelvis|898|Carcinosarcoma|8980/3|Carcinosarcoma
C659, C669|RenalPelvis|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C659, C669|RenalPelvis|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C659, C669|RenalPelvis|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C659, C669|RenalPelvis|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C659, C669|RenalPelvis|950|Neuroblastoma|9500/3|Neuroblastoma
C659, C669|RenalPelvis|950|Neuroblastoma|9501/3|Medulloepithelioma
C659, C669|RenalPelvis|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C659, C669|RenalPelvis|950|Neuroblastoma|9503/3|Neuroepithelioma
C659, C669|RenalPelvis|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C659, C669|RenalPelvis|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C659, C669|RenalPelvis|959|Lymphoma|9590/3|Lymphoma
C659, C669|RenalPelvis|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C659, C669|RenalPelvis|959|Lymphoma|9596/3|CompositeLymphoma
C659, C669|RenalPelvis|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C659, C669|RenalPelvis|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C659, C669|RenalPelvis|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C659, C669|RenalPelvis|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C659, C669|RenalPelvis|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C659, C669|RenalPelvis|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C659, C669|RenalPelvis|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C659, C669|RenalPelvis|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C659, C669|RenalPelvis|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C659, C669|RenalPelvis|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C659, C669|RenalPelvis|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C659, C669|RenalPelvis|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C659, C669|RenalPelvis|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C659, C669|RenalPelvis|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C659, C669|RenalPelvis|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C659, C669|RenalPelvis|967|BCellLymphomas|9673/3|MantleCellLymphoma
C659, C669|RenalPelvis|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C659, C669|RenalPelvis|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C659, C669|RenalPelvis|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C659, C669|RenalPelvis|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C659, C669|RenalPelvis|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C659, C669|RenalPelvis|969|FollicularAdenoma|9690/3|LymphomaFollicular
C659, C669|RenalPelvis|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C659, C669|RenalPelvis|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C659, C669|RenalPelvis|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C659, C669|RenalPelvis|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C659, C669|RenalPelvis|970|TCellLymphoma|9701/3|SezarySyndrome
C659, C669|RenalPelvis|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C659, C669|RenalPelvis|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C659, C669|RenalPelvis|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C659, C669|RenalPelvis|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C659, C669|RenalPelvis|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C659, C669|RenalPelvis|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C659, C669|RenalPelvis|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C659, C669|RenalPelvis|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C659, C669|RenalPelvis|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C659, C669|RenalPelvis|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C659, C669|RenalPelvis|973|Plasmacytoma|9731/3|Plasmacytoma
C659, C669|RenalPelvis|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C659, C669|RenalPelvis|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C659, C669|RenalPelvis|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C659, C669|RenalPelvis|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C659, C669|RenalPelvis|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C659, C669|RenalPelvis|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C659, C669|RenalPelvis|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C659, C669|RenalPelvis|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C659, C669|RenalPelvis|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C659, C669|RenalPelvis|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C659, C669|RenalPelvis|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C659, C669|RenalPelvis|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C659, C669|RenalPelvis|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C659, C669|RenalPelvis|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C659, C669|RenalPelvis|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C659, C669|RenalPelvis|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9812/3|null
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9813/3|null
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9814/3|null
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9817/3|null
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9818/3|null
C659, C669|RenalPelvis|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C659, C669|RenalPelvis|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C659, C669|RenalPelvis|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C659, C669|RenalPelvis|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C659, C669|RenalPelvis|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C659, C669|RenalPelvis|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C659, C669|RenalPelvis|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C659, C669|RenalPelvis|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C670-C679|UrinaryBladder|801|Carcinoma|8010/2|InSituCancer
C670-C679|UrinaryBladder|801|Carcinoma|8010/3|CarcinomaNOSDNE
C670-C679|UrinaryBladder|801|Carcinoma|8011/3|MalignantEpithelioma
C670-C679|UrinaryBladder|801|Carcinoma|8012/3|LargeCellCarcinoma
C670-C679|UrinaryBladder|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C670-C679|UrinaryBladder|801|Carcinoma|8014/3|LargeCellCarcinoma
C670-C679|UrinaryBladder|801|Carcinoma|8015/3|GlassyCellCarcinoma
C670-C679|UrinaryBladder|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C670-C679|UrinaryBladder|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C670-C679|UrinaryBladder|802|Carcinoma|8022/3|PleomorphicCarcinoma
C670-C679|UrinaryBladder|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C670-C679|UrinaryBladder|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C670-C679|UrinaryBladder|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C670-C679|UrinaryBladder|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C670-C679|UrinaryBladder|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C670-C679|UrinaryBladder|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C670-C679|UrinaryBladder|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C670-C679|UrinaryBladder|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C670-C679|UrinaryBladder|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C670-C679|UrinaryBladder|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C670-C679|UrinaryBladder|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C670-C679|UrinaryBladder|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C670-C679|UrinaryBladder|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C670-C679|UrinaryBladder|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C670-C679|UrinaryBladder|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C670-C679|UrinaryBladder|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C670-C679|UrinaryBladder|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C670-C679|UrinaryBladder|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C670-C679|UrinaryBladder|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C670-C679|UrinaryBladder|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C670-C679|UrinaryBladder|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C670-C679|UrinaryBladder|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C670-C679|UrinaryBladder|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C670-C679|UrinaryBladder|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C670-C679|UrinaryBladder|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C670-C679|UrinaryBladder|814|Adenocarcinoma|8140/3|Adenocarcinoma
C670-C679|UrinaryBladder|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C670-C679|UrinaryBladder|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C670-C679|UrinaryBladder|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C670-C679|UrinaryBladder|823|SolidCarcinoma|8230/2|InSituCancer
C670-C679|UrinaryBladder|823|SolidCarcinoma|8230/3|SolidCarcinoma
C670-C679|UrinaryBladder|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C670-C679|UrinaryBladder|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C670-C679|UrinaryBladder|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C670-C679|UrinaryBladder|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C670-C679|UrinaryBladder|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C670-C679|UrinaryBladder|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C670-C679|UrinaryBladder|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C670-C679|UrinaryBladder|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C670-C679|UrinaryBladder|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C670-C679|UrinaryBladder|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C670-C679|UrinaryBladder|849|SignetRingCellCarcinoma|8490/3|SignetRingCellCarcinoma
C670-C679|UrinaryBladder|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C670-C679|UrinaryBladder|857|AdenocarcinomaWithMetaplasia|8576/3|HepatoidAdenocarcinoma
C670-C679|UrinaryBladder|868|Paraganglioma|8680/3|MalignantParaganglioma
C670-C679|UrinaryBladder|880|Sarcoma|8800/3|Sarcoma
C670-C679|UrinaryBladder|880|Sarcoma|8801/3|SpindleCellSarcoma
C670-C679|UrinaryBladder|880|Sarcoma|8802/3|GiantCellSarcoma
C670-C679|UrinaryBladder|880|Sarcoma|8803/3|SmallCellSarcoma
C670-C679|UrinaryBladder|880|Sarcoma|8804/3|SarcomaEpithelioid
C670-C679|UrinaryBladder|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C670-C679|UrinaryBladder|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C670-C679|UrinaryBladder|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C670-C679|UrinaryBladder|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C670-C679|UrinaryBladder|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C670-C679|UrinaryBladder|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C670-C679|UrinaryBladder|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C670-C679|UrinaryBladder|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C670-C679|UrinaryBladder|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C670-C679|UrinaryBladder|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C670-C679|UrinaryBladder|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C670-C679|UrinaryBladder|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C670-C679|UrinaryBladder|889|MyomatousNeoplasm|8895/3|Myosarcoma
C670-C679|UrinaryBladder|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C670-C679|UrinaryBladder|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C670-C679|UrinaryBladder|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C670-C679|UrinaryBladder|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C670-C679|UrinaryBladder|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C670-C679|UrinaryBladder|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C670-C679|UrinaryBladder|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C670-C679|UrinaryBladder|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C670-C679|UrinaryBladder|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C670-C679|UrinaryBladder|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C670-C679|UrinaryBladder|898|Carcinosarcoma|8980/3|Carcinosarcoma
C670-C679|UrinaryBladder|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C670-C679|UrinaryBladder|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C670-C679|UrinaryBladder|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C670-C679|UrinaryBladder|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C670-C679|UrinaryBladder|959|Lymphoma|9590/3|Lymphoma
C670-C679|UrinaryBladder|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C670-C679|UrinaryBladder|959|Lymphoma|9596/3|CompositeLymphoma
C670-C679|UrinaryBladder|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C670-C679|UrinaryBladder|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C670-C679|UrinaryBladder|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C670-C679|UrinaryBladder|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C670-C679|UrinaryBladder|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C670-C679|UrinaryBladder|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C670-C679|UrinaryBladder|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C670-C679|UrinaryBladder|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C670-C679|UrinaryBladder|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C670-C679|UrinaryBladder|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C670-C679|UrinaryBladder|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C670-C679|UrinaryBladder|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C670-C679|UrinaryBladder|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C670-C679|UrinaryBladder|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C670-C679|UrinaryBladder|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C670-C679|UrinaryBladder|967|BCellLymphomas|9673/3|MantleCellLymphoma
C670-C679|UrinaryBladder|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C670-C679|UrinaryBladder|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C670-C679|UrinaryBladder|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C670-C679|UrinaryBladder|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C670-C679|UrinaryBladder|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C670-C679|UrinaryBladder|969|FollicularAdenoma|9690/3|LymphomaFollicular
C670-C679|UrinaryBladder|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C670-C679|UrinaryBladder|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C670-C679|UrinaryBladder|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C670-C679|UrinaryBladder|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C670-C679|UrinaryBladder|970|TCellLymphoma|9701/3|SezarySyndrome
C670-C679|UrinaryBladder|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C670-C679|UrinaryBladder|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C670-C679|UrinaryBladder|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C670-C679|UrinaryBladder|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C670-C679|UrinaryBladder|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C670-C679|UrinaryBladder|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C670-C679|UrinaryBladder|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C670-C679|UrinaryBladder|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C670-C679|UrinaryBladder|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C670-C679|UrinaryBladder|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C670-C679|UrinaryBladder|973|Plasmacytoma|9731/3|Plasmacytoma
C670-C679|UrinaryBladder|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C670-C679|UrinaryBladder|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C670-C679|UrinaryBladder|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C670-C679|UrinaryBladder|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C670-C679|UrinaryBladder|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C670-C679|UrinaryBladder|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C670-C679|UrinaryBladder|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C670-C679|UrinaryBladder|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C670-C679|UrinaryBladder|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C670-C679|UrinaryBladder|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C670-C679|UrinaryBladder|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C670-C679|UrinaryBladder|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C670-C679|UrinaryBladder|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C670-C679|UrinaryBladder|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C670-C679|UrinaryBladder|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C670-C679|UrinaryBladder|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9812/3|null
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9813/3|null
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9814/3|null
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9817/3|null
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9818/3|null
C670-C679|UrinaryBladder|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C670-C679|UrinaryBladder|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C670-C679|UrinaryBladder|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C670-C679|UrinaryBladder|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C670-C679|UrinaryBladder|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C670-C679|UrinaryBladder|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C670-C679|UrinaryBladder|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C670-C679|UrinaryBladder|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C680-C681,C688-C689|GenitourinarySystem|801|Carcinoma|8010/2|InSituCancer
C680-C681,C688-C689|GenitourinarySystem|801|Carcinoma|8010/3|CarcinomaNOSDNE
C680-C681,C688-C689|GenitourinarySystem|801|Carcinoma|8011/3|MalignantEpithelioma
C680-C681,C688-C689|GenitourinarySystem|801|Carcinoma|8012/3|LargeCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C680-C681,C688-C689|GenitourinarySystem|801|Carcinoma|8014/3|LargeCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|801|Carcinoma|8015/3|GlassyCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C680-C681,C688-C689|GenitourinarySystem|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C680-C681,C688-C689|GenitourinarySystem|802|Carcinoma|8022/3|PleomorphicCarcinoma
C680-C681,C688-C689|GenitourinarySystem|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C680-C681,C688-C689|GenitourinarySystem|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C680-C681,C688-C689|GenitourinarySystem|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C680-C681,C688-C689|GenitourinarySystem|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C680-C681,C688-C689|GenitourinarySystem|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C680-C681,C688-C689|GenitourinarySystem|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C680-C681,C688-C689|GenitourinarySystem|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C680-C681,C688-C689|GenitourinarySystem|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C680-C681,C688-C689|GenitourinarySystem|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C680-C681,C688-C689|GenitourinarySystem|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C680-C681,C688-C689|GenitourinarySystem|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C680-C681,C688-C689|GenitourinarySystem|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C680-C681,C688-C689|GenitourinarySystem|814|Adenocarcinoma|8140/3|Adenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C680-C681,C688-C689|GenitourinarySystem|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|823|SolidCarcinoma|8230/2|InSituCancer
C680-C681,C688-C689|GenitourinarySystem|823|SolidCarcinoma|8230/3|SolidCarcinoma
C680-C681,C688-C689|GenitourinarySystem|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C680-C681,C688-C689|GenitourinarySystem|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C680-C681,C688-C689|GenitourinarySystem|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C680-C681,C688-C689|GenitourinarySystem|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C680-C681,C688-C689|GenitourinarySystem|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C680-C681,C688-C689|GenitourinarySystem|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C680-C681,C688-C689|GenitourinarySystem|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C680-C681,C688-C689|GenitourinarySystem|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|838|CarcinomaEndometrioid|8380/3|CarcinomaEndometrioid
C680-C681,C688-C689|GenitourinarySystem|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|848|MucinousAdenocarcinoma|8480/3|MucinousAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|848|MucinousAdenocarcinoma|8481/3|MucinProducingAdenocarcinoma
C680-C681,C688-C689|GenitourinarySystem|856|AdenosquamousCarcinoma|8560/3|AdenosquamousCarcinoma
C680-C681,C688-C689|GenitourinarySystem|856|AdenosquamousCarcinoma|8562/3|EpithelialMyoepithelialCarcinoma
C680-C681,C688-C689|GenitourinarySystem|872|Melanoma|8720/2|Stage0SkinMelanoma
C680-C681,C688-C689|GenitourinarySystem|872|Melanoma|8720/3|Melanoma
C680-C681,C688-C689|GenitourinarySystem|872|Melanoma|8721/3|NodularMelanoma
C680-C681,C688-C689|GenitourinarySystem|872|Melanoma|8722/3|BalloonCellMelanoma
C680-C681,C688-C689|GenitourinarySystem|872|Melanoma|8723/3|RegressingMelanoma
C680-C681,C688-C689|GenitourinarySystem|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C680-C681,C688-C689|GenitourinarySystem|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C680-C681,C688-C689|GenitourinarySystem|874|Nevus|8745/3|DesmoplasticMelanoma
C680-C681,C688-C689|GenitourinarySystem|874|Nevus|8746/3|MucosalLentiginousMelanoma
C680-C681,C688-C689|GenitourinarySystem|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C680-C681,C688-C689|GenitourinarySystem|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C680-C681,C688-C689|GenitourinarySystem|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C680-C681,C688-C689|GenitourinarySystem|880|Sarcoma|8800/3|Sarcoma
C680-C681,C688-C689|GenitourinarySystem|880|Sarcoma|8801/3|SpindleCellSarcoma
C680-C681,C688-C689|GenitourinarySystem|880|Sarcoma|8802/3|GiantCellSarcoma
C680-C681,C688-C689|GenitourinarySystem|880|Sarcoma|8803/3|SmallCellSarcoma
C680-C681,C688-C689|GenitourinarySystem|880|Sarcoma|8804/3|SarcomaEpithelioid
C680-C681,C688-C689|GenitourinarySystem|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C680-C681,C688-C689|GenitourinarySystem|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C680-C681,C688-C689|GenitourinarySystem|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C680-C681,C688-C689|GenitourinarySystem|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C680-C681,C688-C689|GenitourinarySystem|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C680-C681,C688-C689|GenitourinarySystem|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C680-C681,C688-C689|GenitourinarySystem|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C680-C681,C688-C689|GenitourinarySystem|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C680-C681,C688-C689|GenitourinarySystem|885|Liposarcoma|8850/3|Liposarcoma
C680-C681,C688-C689|GenitourinarySystem|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C680-C681,C688-C689|GenitourinarySystem|885|Liposarcoma|8852/3|LiposarcomaMyxoid
C680-C681,C688-C689|GenitourinarySystem|885|Liposarcoma|8853/3|RoundCellLiposarcoma
C680-C681,C688-C689|GenitourinarySystem|885|Liposarcoma|8854/3|PleomorphicLiposarcoma
C680-C681,C688-C689|GenitourinarySystem|885|Liposarcoma|8855/3|Liposarcoma
C680-C681,C688-C689|GenitourinarySystem|885|Liposarcoma|8857/3|FibroblasticLiposarcoma
C680-C681,C688-C689|GenitourinarySystem|885|Liposarcoma|8858/3|DedifferentiatedLiposarcoma
C680-C681,C688-C689|GenitourinarySystem|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|889|MyomatousNeoplasm|8895/3|Myosarcoma
C680-C681,C688-C689|GenitourinarySystem|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C680-C681,C688-C689|GenitourinarySystem|895|MixedTumorMullerian|8950/3|MixedTumorMullerian
C680-C681,C688-C689|GenitourinarySystem|895|MixedTumorMullerian|8951/3|MesodermalMixedTumor
C680-C681,C688-C689|GenitourinarySystem|896|Nephroblastoma|8964/3|ClearCellSarcomaOfTheKidney
C680-C681,C688-C689|GenitourinarySystem|898|Carcinosarcoma|8980/3|Carcinosarcoma
C680-C681,C688-C689|GenitourinarySystem|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C680-C681,C688-C689|GenitourinarySystem|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C680-C681,C688-C689|GenitourinarySystem|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C680-C681,C688-C689|GenitourinarySystem|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C680-C681,C688-C689|GenitourinarySystem|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C680-C681,C688-C689|GenitourinarySystem|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C680-C681,C688-C689|GenitourinarySystem|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C680-C681,C688-C689|GenitourinarySystem|908|Teratoma|9080/3|ImmatureTeratoma
C680-C681,C688-C689|GenitourinarySystem|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C680-C681,C688-C689|GenitourinarySystem|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C680-C681,C688-C689|GenitourinarySystem|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C680-C681,C688-C689|GenitourinarySystem|908|Teratoma|9084/3|Teratoma
C680-C681,C688-C689|GenitourinarySystem|908|Teratoma|9085/3|MixedGermCellTumor
C680-C681,C688-C689|GenitourinarySystem|911|Mesonephroma|9110/3|Mesonephroma
C680-C681,C688-C689|GenitourinarySystem|950|Neuroblastoma|9500/3|Neuroblastoma
C680-C681,C688-C689|GenitourinarySystem|950|Neuroblastoma|9501/3|Medulloepithelioma
C680-C681,C688-C689|GenitourinarySystem|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C680-C681,C688-C689|GenitourinarySystem|950|Neuroblastoma|9503/3|Neuroepithelioma
C680-C681,C688-C689|GenitourinarySystem|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C680-C681,C688-C689|GenitourinarySystem|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C680-C681,C688-C689|GenitourinarySystem|959|Lymphoma|9590/3|Lymphoma
C680-C681,C688-C689|GenitourinarySystem|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C680-C681,C688-C689|GenitourinarySystem|959|Lymphoma|9596/3|CompositeLymphoma
C680-C681,C688-C689|GenitourinarySystem|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C680-C681,C688-C689|GenitourinarySystem|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C680-C681,C688-C689|GenitourinarySystem|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C680-C681,C688-C689|GenitourinarySystem|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C680-C681,C688-C689|GenitourinarySystem|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C680-C681,C688-C689|GenitourinarySystem|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C680-C681,C688-C689|GenitourinarySystem|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C680-C681,C688-C689|GenitourinarySystem|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C680-C681,C688-C689|GenitourinarySystem|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C680-C681,C688-C689|GenitourinarySystem|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C680-C681,C688-C689|GenitourinarySystem|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C680-C681,C688-C689|GenitourinarySystem|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C680-C681,C688-C689|GenitourinarySystem|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C680-C681,C688-C689|GenitourinarySystem|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C680-C681,C688-C689|GenitourinarySystem|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C680-C681,C688-C689|GenitourinarySystem|967|BCellLymphomas|9673/3|MantleCellLymphoma
C680-C681,C688-C689|GenitourinarySystem|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C680-C681,C688-C689|GenitourinarySystem|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C680-C681,C688-C689|GenitourinarySystem|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C680-C681,C688-C689|GenitourinarySystem|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C680-C681,C688-C689|GenitourinarySystem|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C680-C681,C688-C689|GenitourinarySystem|969|FollicularAdenoma|9690/3|LymphomaFollicular
C680-C681,C688-C689|GenitourinarySystem|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C680-C681,C688-C689|GenitourinarySystem|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C680-C681,C688-C689|GenitourinarySystem|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C680-C681,C688-C689|GenitourinarySystem|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C680-C681,C688-C689|GenitourinarySystem|970|TCellLymphoma|9701/3|SezarySyndrome
C680-C681,C688-C689|GenitourinarySystem|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C680-C681,C688-C689|GenitourinarySystem|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C680-C681,C688-C689|GenitourinarySystem|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C680-C681,C688-C689|GenitourinarySystem|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C680-C681,C688-C689|GenitourinarySystem|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C680-C681,C688-C689|GenitourinarySystem|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C680-C681,C688-C689|GenitourinarySystem|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C680-C681,C688-C689|GenitourinarySystem|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C680-C681,C688-C689|GenitourinarySystem|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C680-C681,C688-C689|GenitourinarySystem|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C680-C681,C688-C689|GenitourinarySystem|973|Plasmacytoma|9731/3|Plasmacytoma
C680-C681,C688-C689|GenitourinarySystem|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C680-C681,C688-C689|GenitourinarySystem|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C680-C681,C688-C689|GenitourinarySystem|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C680-C681,C688-C689|GenitourinarySystem|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C680-C681,C688-C689|GenitourinarySystem|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C680-C681,C688-C689|GenitourinarySystem|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C680-C681,C688-C689|GenitourinarySystem|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C680-C681,C688-C689|GenitourinarySystem|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C680-C681,C688-C689|GenitourinarySystem|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C680-C681,C688-C689|GenitourinarySystem|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C680-C681,C688-C689|GenitourinarySystem|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C680-C681,C688-C689|GenitourinarySystem|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C680-C681,C688-C689|GenitourinarySystem|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C680-C681,C688-C689|GenitourinarySystem|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C680-C681,C688-C689|GenitourinarySystem|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C680-C681,C688-C689|GenitourinarySystem|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9812/3|null
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9813/3|null
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9814/3|null
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9817/3|null
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9818/3|null
C680-C681,C688-C689|GenitourinarySystem|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C680-C681,C688-C689|GenitourinarySystem|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C680-C681,C688-C689|GenitourinarySystem|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C680-C681,C688-C689|GenitourinarySystem|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C680-C681,C688-C689|GenitourinarySystem|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C680-C681,C688-C689|GenitourinarySystem|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C680-C681,C688-C689|GenitourinarySystem|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C680-C681,C688-C689|GenitourinarySystem|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C690-C691, C693, C695-C698|LacrimalGland|801|Carcinoma|8010/2|InSituCancer
C690-C691, C693, C695-C698|LacrimalGland|801|Carcinoma|8010/3|CarcinomaNOSDNE
C690-C691, C693, C695-C698|LacrimalGland|801|Carcinoma|8011/3|MalignantEpithelioma
C690-C691, C693, C695-C698|LacrimalGland|801|Carcinoma|8012/3|LargeCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|801|Carcinoma|8014/3|LargeCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|801|Carcinoma|8015/3|GlassyCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C690-C691, C693, C695-C698|LacrimalGland|802|Carcinoma|8022/3|PleomorphicCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C690-C691, C693, C695-C698|LacrimalGland|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C690-C691, C693, C695-C698|LacrimalGland|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C690-C691, C693, C695-C698|LacrimalGland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C690-C691, C693, C695-C698|LacrimalGland|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C690-C691, C693, C695-C698|LacrimalGland|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C690-C691, C693, C695-C698|LacrimalGland|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C690-C691, C693, C695-C698|LacrimalGland|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C690-C691, C693, C695-C698|LacrimalGland|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C690-C691, C693, C695-C698|LacrimalGland|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C690-C691, C693, C695-C698|LacrimalGland|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C690-C691, C693, C695-C698|LacrimalGland|872|Melanoma|8720/2|Stage0SkinMelanoma
C690-C691, C693, C695-C698|LacrimalGland|872|Melanoma|8720/3|Melanoma
C690-C691, C693, C695-C698|LacrimalGland|872|Melanoma|8721/3|NodularMelanoma
C690-C691, C693, C695-C698|LacrimalGland|872|Melanoma|8722/3|BalloonCellMelanoma
C690-C691, C693, C695-C698|LacrimalGland|872|Melanoma|8723/3|RegressingMelanoma
C690-C691, C693, C695-C698|LacrimalGland|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C690-C691, C693, C695-C698|LacrimalGland|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C690-C691, C693, C695-C698|LacrimalGland|874|Nevus|8745/3|DesmoplasticMelanoma
C690-C691, C693, C695-C698|LacrimalGland|874|Nevus|8746/3|MucosalLentiginousMelanoma
C690-C691, C693, C695-C698|LacrimalGland|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C690-C691, C693, C695-C698|LacrimalGland|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C690-C691, C693, C695-C698|LacrimalGland|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C690-C691, C693, C695-C698|LacrimalGland|877|EpithelioidCellMelanoma|8773/3|TypeASpindleCellMelanoma
C690-C691, C693, C695-C698|LacrimalGland|877|EpithelioidCellMelanoma|8774/3|TypeBSpindleCellMelanoma
C690-C691, C693, C695-C698|LacrimalGland|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C690-C691, C693, C695-C698|LacrimalGland|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C690-C691, C693, C695-C698|LacrimalGland|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C690-C691, C693, C695-C698|LacrimalGland|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C690-C691, C693, C695-C698|LacrimalGland|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C690-C691, C693, C695-C698|LacrimalGland|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C690-C691, C693, C695-C698|LacrimalGland|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|889|MyomatousNeoplasm|8895/3|Myosarcoma
C690-C691, C693, C695-C698|LacrimalGland|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C690-C691, C693, C695-C698|LacrimalGland|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C690-C691, C693, C695-C698|LacrimalGland|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C690-C691, C693, C695-C698|LacrimalGland|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C690-C691, C693, C695-C698|LacrimalGland|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C690-C691, C693, C695-C698|LacrimalGland|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C690-C691, C693, C695-C698|LacrimalGland|959|Lymphoma|9590/3|Lymphoma
C690-C691, C693, C695-C698|LacrimalGland|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C690-C691, C693, C695-C698|LacrimalGland|959|Lymphoma|9596/3|CompositeLymphoma
C690-C691, C693, C695-C698|LacrimalGland|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C690-C691, C693, C695-C698|LacrimalGland|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C690-C691, C693, C695-C698|LacrimalGland|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C690-C691, C693, C695-C698|LacrimalGland|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C690-C691, C693, C695-C698|LacrimalGland|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C690-C691, C693, C695-C698|LacrimalGland|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C690-C691, C693, C695-C698|LacrimalGland|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C690-C691, C693, C695-C698|LacrimalGland|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C690-C691, C693, C695-C698|LacrimalGland|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C690-C691, C693, C695-C698|LacrimalGland|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C690-C691, C693, C695-C698|LacrimalGland|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C690-C691, C693, C695-C698|LacrimalGland|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C690-C691, C693, C695-C698|LacrimalGland|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C690-C691, C693, C695-C698|LacrimalGland|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C690-C691, C693, C695-C698|LacrimalGland|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C690-C691, C693, C695-C698|LacrimalGland|967|BCellLymphomas|9673/3|MantleCellLymphoma
C690-C691, C693, C695-C698|LacrimalGland|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C690-C691, C693, C695-C698|LacrimalGland|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C690-C691, C693, C695-C698|LacrimalGland|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C690-C691, C693, C695-C698|LacrimalGland|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C690-C691, C693, C695-C698|LacrimalGland|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C690-C691, C693, C695-C698|LacrimalGland|969|FollicularAdenoma|9690/3|LymphomaFollicular
C690-C691, C693, C695-C698|LacrimalGland|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C690-C691, C693, C695-C698|LacrimalGland|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C690-C691, C693, C695-C698|LacrimalGland|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C690-C691, C693, C695-C698|LacrimalGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C690-C691, C693, C695-C698|LacrimalGland|970|TCellLymphoma|9701/3|SezarySyndrome
C690-C691, C693, C695-C698|LacrimalGland|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C690-C691, C693, C695-C698|LacrimalGland|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C690-C691, C693, C695-C698|LacrimalGland|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C690-C691, C693, C695-C698|LacrimalGland|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C690-C691, C693, C695-C698|LacrimalGland|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C690-C691, C693, C695-C698|LacrimalGland|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C690-C691, C693, C695-C698|LacrimalGland|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C690-C691, C693, C695-C698|LacrimalGland|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C690-C691, C693, C695-C698|LacrimalGland|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C690-C691, C693, C695-C698|LacrimalGland|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C690-C691, C693, C695-C698|LacrimalGland|973|Plasmacytoma|9731/3|Plasmacytoma
C690-C691, C693, C695-C698|LacrimalGland|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C690-C691, C693, C695-C698|LacrimalGland|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C690-C691, C693, C695-C698|LacrimalGland|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C690-C691, C693, C695-C698|LacrimalGland|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C690-C691, C693, C695-C698|LacrimalGland|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C690-C691, C693, C695-C698|LacrimalGland|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C690-C691, C693, C695-C698|LacrimalGland|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C690-C691, C693, C695-C698|LacrimalGland|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C690-C691, C693, C695-C698|LacrimalGland|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C690-C691, C693, C695-C698|LacrimalGland|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C690-C691, C693, C695-C698|LacrimalGland|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C690-C691, C693, C695-C698|LacrimalGland|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C690-C691, C693, C695-C698|LacrimalGland|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C690-C691, C693, C695-C698|LacrimalGland|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C690-C691, C693, C695-C698|LacrimalGland|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C690-C691, C693, C695-C698|LacrimalGland|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9812/3|null
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9813/3|null
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9814/3|null
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9817/3|null
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9818/3|null
C690-C691, C693, C695-C698|LacrimalGland|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C690-C691, C693, C695-C698|LacrimalGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C690-C691, C693, C695-C698|LacrimalGland|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C690-C691, C693, C695-C698|LacrimalGland|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C690-C691, C693, C695-C698|LacrimalGland|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C690-C691, C693, C695-C698|LacrimalGland|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C690-C691, C693, C695-C698|LacrimalGland|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C690-C691, C693, C695-C698|LacrimalGland|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C692|Retina|801|Carcinoma|8010/2|InSituCancer
C692|Retina|801|Carcinoma|8010/3|CarcinomaNOSDNE
C692|Retina|801|Carcinoma|8011/3|MalignantEpithelioma
C692|Retina|801|Carcinoma|8012/3|LargeCellCarcinoma
C692|Retina|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C692|Retina|801|Carcinoma|8014/3|LargeCellCarcinoma
C692|Retina|801|Carcinoma|8015/3|GlassyCellCarcinoma
C692|Retina|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C692|Retina|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C692|Retina|802|Carcinoma|8022/3|PleomorphicCarcinoma
C692|Retina|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C692|Retina|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C692|Retina|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C692|Retina|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C692|Retina|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C692|Retina|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C692|Retina|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C692|Retina|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C692|Retina|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C692|Retina|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C692|Retina|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C692|Retina|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C692|Retina|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C692|Retina|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C692|Retina|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C692|Retina|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C692|Retina|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C692|Retina|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C692|Retina|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C692|Retina|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C692|Retina|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C692|Retina|814|Adenocarcinoma|8140/3|Adenocarcinoma
C692|Retina|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C692|Retina|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C692|Retina|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C692|Retina|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C692|Retina|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C692|Retina|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C692|Retina|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C692|Retina|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C692|Retina|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C692|Retina|872|Melanoma|8720/2|Stage0SkinMelanoma
C692|Retina|872|Melanoma|8720/3|Melanoma
C692|Retina|872|Melanoma|8721/3|NodularMelanoma
C692|Retina|872|Melanoma|8722/3|BalloonCellMelanoma
C692|Retina|872|Melanoma|8723/3|RegressingMelanoma
C692|Retina|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C692|Retina|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C692|Retina|874|Nevus|8745/3|DesmoplasticMelanoma
C692|Retina|874|Nevus|8746/3|MucosalLentiginousMelanoma
C692|Retina|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C692|Retina|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C692|Retina|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C692|Retina|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C692|Retina|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C692|Retina|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C692|Retina|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C692|Retina|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C692|Retina|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C692|Retina|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C692|Retina|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C692|Retina|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C692|Retina|889|MyomatousNeoplasm|8895/3|Myosarcoma
C692|Retina|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C692|Retina|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C692|Retina|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C692|Retina|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C692|Retina|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C692|Retina|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C692|Retina|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C692|Retina|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C692|Retina|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C692|Retina|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C692|Retina|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C692|Retina|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C692|Retina|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C692|Retina|951|Retinoblastoma|9510/3|Retinoblastoma
C692|Retina|951|Retinoblastoma|9511/3|DifferentiatedRetinoblastoma
C692|Retina|951|Retinoblastoma|9512/3|UndifferentiatedRetinoblastoma
C692|Retina|951|Retinoblastoma|9513/3|DiffuseRetinoblastoma
C692|Retina|959|Lymphoma|9590/3|Lymphoma
C692|Retina|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C692|Retina|959|Lymphoma|9596/3|CompositeLymphoma
C692|Retina|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C692|Retina|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C692|Retina|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C692|Retina|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C692|Retina|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C692|Retina|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C692|Retina|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C692|Retina|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C692|Retina|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C692|Retina|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C692|Retina|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C692|Retina|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C692|Retina|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C692|Retina|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C692|Retina|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C692|Retina|967|BCellLymphomas|9673/3|MantleCellLymphoma
C692|Retina|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C692|Retina|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C692|Retina|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C692|Retina|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C692|Retina|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C692|Retina|969|FollicularAdenoma|9690/3|LymphomaFollicular
C692|Retina|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C692|Retina|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C692|Retina|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C692|Retina|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C692|Retina|970|TCellLymphoma|9701/3|SezarySyndrome
C692|Retina|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C692|Retina|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C692|Retina|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C692|Retina|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C692|Retina|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C692|Retina|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C692|Retina|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C692|Retina|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C692|Retina|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C692|Retina|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C692|Retina|973|Plasmacytoma|9731/3|Plasmacytoma
C692|Retina|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C692|Retina|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C692|Retina|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C692|Retina|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C692|Retina|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C692|Retina|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C692|Retina|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C692|Retina|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C692|Retina|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C692|Retina|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C692|Retina|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C692|Retina|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C692|Retina|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C692|Retina|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C692|Retina|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C692|Retina|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C692|Retina|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C692|Retina|981|PrecursorLymphoidNeoplasm|9812/3|null
C692|Retina|981|PrecursorLymphoidNeoplasm|9813/3|null
C692|Retina|981|PrecursorLymphoidNeoplasm|9814/3|null
C692|Retina|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C692|Retina|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C692|Retina|981|PrecursorLymphoidNeoplasm|9817/3|null
C692|Retina|981|PrecursorLymphoidNeoplasm|9818/3|null
C692|Retina|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C692|Retina|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C692|Retina|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C692|Retina|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C692|Retina|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C692|Retina|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C692|Retina|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C692|Retina|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C694|Eye|801|Carcinoma|8010/2|InSituCancer
C694|Eye|801|Carcinoma|8010/3|CarcinomaNOSDNE
C694|Eye|801|Carcinoma|8011/3|MalignantEpithelioma
C694|Eye|801|Carcinoma|8012/3|LargeCellCarcinoma
C694|Eye|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C694|Eye|801|Carcinoma|8014/3|LargeCellCarcinoma
C694|Eye|801|Carcinoma|8015/3|GlassyCellCarcinoma
C694|Eye|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C694|Eye|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C694|Eye|802|Carcinoma|8022/3|PleomorphicCarcinoma
C694|Eye|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C694|Eye|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C694|Eye|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C694|Eye|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C694|Eye|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C694|Eye|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C694|Eye|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C694|Eye|808|LymphoepithelialCarcinoma|8081/2|BowenDisease
C694|Eye|808|LymphoepithelialCarcinoma|8082/3|LymphoepithelialCarcinoma
C694|Eye|808|LymphoepithelialCarcinoma|8083/3|BasaloidSquamousCellCarcinoma
C694|Eye|808|LymphoepithelialCarcinoma|8084/3|ClearCellSquamousCellSkinCarcinoma
C694|Eye|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C694|Eye|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C694|Eye|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C694|Eye|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C694|Eye|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C694|Eye|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C694|Eye|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C694|Eye|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C694|Eye|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C694|Eye|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C694|Eye|814|Adenocarcinoma|8140/3|Adenocarcinoma
C694|Eye|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C694|Eye|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C694|Eye|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C694|Eye|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C694|Eye|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C694|Eye|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C694|Eye|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C694|Eye|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C694|Eye|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C694|Eye|872|Melanoma|8720/2|Stage0SkinMelanoma
C694|Eye|872|Melanoma|8720/3|Melanoma
C694|Eye|872|Melanoma|8721/3|NodularMelanoma
C694|Eye|872|Melanoma|8722/3|BalloonCellMelanoma
C694|Eye|872|Melanoma|8723/3|RegressingMelanoma
C694|Eye|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C694|Eye|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C694|Eye|874|Nevus|8745/3|DesmoplasticMelanoma
C694|Eye|874|Nevus|8746/3|MucosalLentiginousMelanoma
C694|Eye|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C694|Eye|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C694|Eye|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C694|Eye|877|EpithelioidCellMelanoma|8773/3|TypeASpindleCellMelanoma
C694|Eye|877|EpithelioidCellMelanoma|8774/3|TypeBSpindleCellMelanoma
C694|Eye|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C694|Eye|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C694|Eye|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C694|Eye|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C694|Eye|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C694|Eye|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C694|Eye|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C694|Eye|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C694|Eye|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C694|Eye|889|MyomatousNeoplasm|8895/3|Myosarcoma
C694|Eye|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C694|Eye|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C694|Eye|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C694|Eye|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C694|Eye|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C694|Eye|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C694|Eye|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C694|Eye|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C694|Eye|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C694|Eye|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C694|Eye|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C694|Eye|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C694|Eye|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C694|Eye|959|Lymphoma|9590/3|Lymphoma
C694|Eye|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C694|Eye|959|Lymphoma|9596/3|CompositeLymphoma
C694|Eye|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C694|Eye|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C694|Eye|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C694|Eye|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C694|Eye|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C694|Eye|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C694|Eye|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C694|Eye|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C694|Eye|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C694|Eye|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C694|Eye|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C694|Eye|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C694|Eye|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C694|Eye|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C694|Eye|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C694|Eye|967|BCellLymphomas|9673/3|MantleCellLymphoma
C694|Eye|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C694|Eye|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C694|Eye|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C694|Eye|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C694|Eye|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C694|Eye|969|FollicularAdenoma|9690/3|LymphomaFollicular
C694|Eye|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C694|Eye|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C694|Eye|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C694|Eye|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C694|Eye|970|TCellLymphoma|9701/3|SezarySyndrome
C694|Eye|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C694|Eye|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C694|Eye|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C694|Eye|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C694|Eye|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C694|Eye|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C694|Eye|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C694|Eye|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C694|Eye|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C694|Eye|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C694|Eye|973|Plasmacytoma|9731/3|Plasmacytoma
C694|Eye|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C694|Eye|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C694|Eye|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C694|Eye|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C694|Eye|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C694|Eye|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C694|Eye|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C694|Eye|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C694|Eye|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C694|Eye|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C694|Eye|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C694|Eye|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C694|Eye|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C694|Eye|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C694|Eye|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C694|Eye|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C694|Eye|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C694|Eye|981|PrecursorLymphoidNeoplasm|9812/3|null
C694|Eye|981|PrecursorLymphoidNeoplasm|9813/3|null
C694|Eye|981|PrecursorLymphoidNeoplasm|9814/3|null
C694|Eye|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C694|Eye|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C694|Eye|981|PrecursorLymphoidNeoplasm|9817/3|null
C694|Eye|981|PrecursorLymphoidNeoplasm|9818/3|null
C694|Eye|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C694|Eye|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C694|Eye|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C694|Eye|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C694|Eye|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C694|Eye|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C694|Eye|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C694|Eye|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C699|Eye|801|Carcinoma|8010/2|InSituCancer
C699|Eye|801|Carcinoma|8010/3|CarcinomaNOSDNE
C699|Eye|801|Carcinoma|8011/3|MalignantEpithelioma
C699|Eye|801|Carcinoma|8012/3|LargeCellCarcinoma
C699|Eye|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C699|Eye|801|Carcinoma|8014/3|LargeCellCarcinoma
C699|Eye|801|Carcinoma|8015/3|GlassyCellCarcinoma
C699|Eye|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C699|Eye|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C699|Eye|802|Carcinoma|8022/3|PleomorphicCarcinoma
C699|Eye|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C699|Eye|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C699|Eye|805|PapillaryCarcinoma|8051/3|VerrucousCarcinoma
C699|Eye|805|PapillaryCarcinoma|8052/2|PapillarySquamousCellCarcinoma
C699|Eye|805|PapillaryCarcinoma|8052/3|PapillarySquamousCellCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C699|Eye|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C699|Eye|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C699|Eye|812|TransitionalCellCarcinoma|8120/2|Stage0TransitionalCellCarcinoma
C699|Eye|812|TransitionalCellCarcinoma|8120/3|TransitionalCellCarcinoma
C699|Eye|812|TransitionalCellCarcinoma|8121/3|SchneiderianCarcinoma
C699|Eye|812|TransitionalCellCarcinoma|8122/3|SarcomatoidCarcinoma
C699|Eye|812|TransitionalCellCarcinoma|8123/3|BasaloidCarcinoma
C699|Eye|812|TransitionalCellCarcinoma|8124/3|AnalCanalCloacogenicCarcinoma
C699|Eye|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C699|Eye|813|PapillaryTransitionalCellCarcinoma|8130/2|PapillaryTransitionalCellCarcinoma
C699|Eye|813|TransitionalCellCarcinoma|8131/3|TransitionalCellCarcinoma
C699|Eye|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C699|Eye|814|Adenocarcinoma|8140/3|Adenocarcinoma
C699|Eye|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C699|Eye|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C699|Eye|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C699|Eye|820|CribriformCarcinoma|8200/3|AdenoidCysticCarcinoma
C699|Eye|820|CribriformCarcinoma|8201/2|CribriformCarcinomaInSitu
C699|Eye|820|CribriformCarcinoma|8201/3|CribriformCarcinoma
C699|Eye|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C699|Eye|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C699|Eye|843|MucoepidermoidCarcinoma|8430/3|MucoepidermoidCarcinoma
C699|Eye|872|Melanoma|8720/2|Stage0SkinMelanoma
C699|Eye|872|Melanoma|8720/3|Melanoma
C699|Eye|872|Melanoma|8721/3|NodularMelanoma
C699|Eye|872|Melanoma|8722/3|BalloonCellMelanoma
C699|Eye|872|Melanoma|8723/3|RegressingMelanoma
C699|Eye|873|MelanomaAmelanotic|8730/3|MelanomaAmelanotic
C699|Eye|874|Nevus|8743/3|SuperficialSpreadingMelanoma
C699|Eye|874|Nevus|8745/3|DesmoplasticMelanoma
C699|Eye|874|Nevus|8746/3|MucosalLentiginousMelanoma
C699|Eye|877|EpithelioidCellMelanoma|8770/3|SpindleCellMelanoma
C699|Eye|877|EpithelioidCellMelanoma|8771/3|EpithelioidCellMelanoma
C699|Eye|877|EpithelioidCellMelanoma|8772/3|SpindleCellMelanoma
C699|Eye|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C699|Eye|881|FibromatousNeoplasm|8811/3|Myxofibrosarcoma
C699|Eye|881|FibromatousNeoplasm|8813/3|FascialFibrosarcoma
C699|Eye|881|FibromatousNeoplasm|8814/3|InfantileFibrosarcoma
C699|Eye|881|FibromatousNeoplasm|8815/3|MalignantSolitaryFibrousTumor
C699|Eye|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C699|Eye|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C699|Eye|889|MyomatousNeoplasm|8891/3|EpithelioidLeiomyosarcoma
C699|Eye|889|MyomatousNeoplasm|8894/3|Angiomyosarcoma
C699|Eye|889|MyomatousNeoplasm|8895/3|Myosarcoma
C699|Eye|889|MyomatousNeoplasm|8896/3|MyxoidLeiomyosarcoma
C699|Eye|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C699|Eye|890|Rhabdomyosarcoma|8901/3|PleomorphicRhabdomyosarcoma
C699|Eye|890|Rhabdomyosarcoma|8902/3|MixedTypeRhabdomyosarcoma
C699|Eye|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C699|Eye|891|EmbryonalRhabdomyosarcoma|8912/3|SpindleCellRhabdomyosarcoma
C699|Eye|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C699|Eye|892|AlveolarRhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C699|Eye|894|MalignantMixedTumor|8940/3|MalignantMixedTumor
C699|Eye|894|MalignantMixedTumor|8941/3|CarcinomaExPleomorphicAdenoma
C699|Eye|899|MalignantMesenchymoma|8990/3|MalignantMesenchymoma
C699|Eye|899|MalignantMesenchymoma|8991/3|UndifferentiatedEmbryonalSarcoma
C699|Eye|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C699|Eye|951|Retinoblastoma|9510/3|Retinoblastoma
C699|Eye|951|Retinoblastoma|9511/3|DifferentiatedRetinoblastoma
C699|Eye|951|Retinoblastoma|9512/3|UndifferentiatedRetinoblastoma
C699|Eye|951|Retinoblastoma|9513/3|DiffuseRetinoblastoma
C699|Eye|959|Lymphoma|9590/3|Lymphoma
C699|Eye|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C699|Eye|959|Lymphoma|9596/3|CompositeLymphoma
C699|Eye|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C699|Eye|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C699|Eye|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C699|Eye|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C699|Eye|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C699|Eye|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C699|Eye|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C699|Eye|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C699|Eye|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C699|Eye|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C699|Eye|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C699|Eye|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C699|Eye|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C699|Eye|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C699|Eye|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C699|Eye|967|BCellLymphomas|9673/3|MantleCellLymphoma
C699|Eye|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C699|Eye|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C699|Eye|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C699|Eye|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C699|Eye|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C699|Eye|969|FollicularAdenoma|9690/3|LymphomaFollicular
C699|Eye|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C699|Eye|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C699|Eye|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C699|Eye|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C699|Eye|970|TCellLymphoma|9701/3|SezarySyndrome
C699|Eye|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C699|Eye|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C699|Eye|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C699|Eye|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C699|Eye|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C699|Eye|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C699|Eye|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C699|Eye|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C699|Eye|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C699|Eye|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C699|Eye|973|Plasmacytoma|9731/3|Plasmacytoma
C699|Eye|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C699|Eye|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C699|Eye|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C699|Eye|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C699|Eye|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C699|Eye|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C699|Eye|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C699|Eye|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C699|Eye|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C699|Eye|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C699|Eye|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C699|Eye|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C699|Eye|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C699|Eye|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C699|Eye|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C699|Eye|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C699|Eye|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C699|Eye|981|PrecursorLymphoidNeoplasm|9812/3|null
C699|Eye|981|PrecursorLymphoidNeoplasm|9813/3|null
C699|Eye|981|PrecursorLymphoidNeoplasm|9814/3|null
C699|Eye|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C699|Eye|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C699|Eye|981|PrecursorLymphoidNeoplasm|9817/3|null
C699|Eye|981|PrecursorLymphoidNeoplasm|9818/3|null
C699|Eye|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C699|Eye|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C699|Eye|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C699|Eye|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C699|Eye|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C699|Eye|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C699|Eye|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C699|Eye|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C700-C701,C709|Meninges|872|Melanoma|8720/3|Melanoma
C700-C701,C709|Meninges|872|Melanoma|8728/0|MeningealMelanocytosis
C700-C701,C709|Meninges|872|Melanoma|8728/1|MeningealMelanocytoma
C700-C701,C709|Meninges|872|Melanoma|8728/3|MeningealMelanomatosis
C700-C701,C709|Meninges|880|Sarcoma|8800/0|BenignSoftTissueNeoplasm
C700-C701,C709|Meninges|880|Sarcoma|8800/3|Sarcoma
C700-C701,C709|Meninges|880|Sarcoma|8801/3|SpindleCellSarcoma
C700-C701,C709|Meninges|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C700-C701,C709|Meninges|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C700-C701,C709|Meninges|881|FibromatousNeoplasm|8810/0|Fibroma
C700-C701,C709|Meninges|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C700-C701,C709|Meninges|881|FibromatousNeoplasm|8815/0|SolitaryFibrousTumor
C700-C701,C709|Meninges|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C700-C701,C709|Meninges|885|Liposarcoma|8850/0|Lipoma
C700-C701,C709|Meninges|885|Liposarcoma|8851/0|Fibrolipoma
C700-C701,C709|Meninges|886|Angiolipoma|8861/0|Angiolipoma
C700-C701,C709|Meninges|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C700-C701,C709|Meninges|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C700-C701,C709|Meninges|908|Teratoma|9080/0|MatureTeratoma
C700-C701,C709|Meninges|908|Teratoma|9080/1|Teratoma
C700-C701,C709|Meninges|908|Teratoma|9080/3|ImmatureTeratoma
C700-C701,C709|Meninges|908|Teratoma|9084/0|DermoidCyst
C700-C701,C709|Meninges|908|Teratoma|9084/3|Teratoma
C700-C701,C709|Meninges|912|NeoplasmsVascularTissue|9120/0|Hemangioma
C700-C701,C709|Meninges|912|NeoplasmsVascularTissue|9121/0|HemangiomaCavernous
C700-C701,C709|Meninges|915|Hemangiopericytoma|9150/0|BenignHemangiopericytoma
C700-C701,C709|Meninges|915|Hemangiopericytoma|9150/1|Hemangiopericytoma
C700-C701,C709|Meninges|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C700-C701,C709|Meninges|916|Hemangioblastoma|9161/1|Hemangioblastoma
C700-C701,C709|Meninges|924|OsseousAndChondromatousNeoplasms|9240/3|MesenchymalChondrosarcoma
C700-C701,C709|Meninges|953|Meningioma|9530/0|Meningioma
C700-C701,C709|Meninges|953|Meningioma|9530/1|Meningiomatosis
C700-C701,C709|Meninges|953|Meningioma|9530/3|GradeIIIMeningioma
C700-C701,C709|Meninges|953|Meningioma|9531/0|MeningothelialMeningioma
C700-C701,C709|Meninges|953|Meningioma|9532/0|FibrousMeningioma
C700-C701,C709|Meninges|953|Meningioma|9533/0|PsammomatousMeningioma
C700-C701,C709|Meninges|953|Meningioma|9534/0|AngiomatousMeningioma
C700-C701,C709|Meninges|953|Meningioma|9537/0|TransitionalMeningioma
C700-C701,C709|Meninges|953|Meningioma|9538/1|ClearCellMeningioma
C700-C701,C709|Meninges|953|Meningioma|9538/3|PapillaryMeningioma
C700-C701,C709|Meninges|953|Meningioma|9539/1|AtypicalMeningioma
C700-C701,C709|Meninges|953|Meningioma|9539/3|MeningealSarcomatosis
C700-C701,C709|Meninges|959|Lymphoma|9590/3|Lymphoma
C700-C701,C709|Meninges|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C700-C701,C709|Meninges|959|Lymphoma|9596/3|CompositeLymphoma
C700-C701,C709|Meninges|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C700-C701,C709|Meninges|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C700-C701,C709|Meninges|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C700-C701,C709|Meninges|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C700-C701,C709|Meninges|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C700-C701,C709|Meninges|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C700-C701,C709|Meninges|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C700-C701,C709|Meninges|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C700-C701,C709|Meninges|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C700-C701,C709|Meninges|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C700-C701,C709|Meninges|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C700-C701,C709|Meninges|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C700-C701,C709|Meninges|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C700-C701,C709|Meninges|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C700-C701,C709|Meninges|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C700-C701,C709|Meninges|967|BCellLymphomas|9673/3|MantleCellLymphoma
C700-C701,C709|Meninges|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C700-C701,C709|Meninges|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C700-C701,C709|Meninges|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C700-C701,C709|Meninges|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C700-C701,C709|Meninges|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C700-C701,C709|Meninges|969|FollicularAdenoma|9690/3|LymphomaFollicular
C700-C701,C709|Meninges|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C700-C701,C709|Meninges|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C700-C701,C709|Meninges|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C700-C701,C709|Meninges|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C700-C701,C709|Meninges|970|TCellLymphoma|9701/3|SezarySyndrome
C700-C701,C709|Meninges|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C700-C701,C709|Meninges|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C700-C701,C709|Meninges|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C700-C701,C709|Meninges|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C700-C701,C709|Meninges|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C700-C701,C709|Meninges|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C700-C701,C709|Meninges|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C700-C701,C709|Meninges|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C700-C701,C709|Meninges|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C700-C701,C709|Meninges|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C700-C701,C709|Meninges|973|Plasmacytoma|9731/3|Plasmacytoma
C700-C701,C709|Meninges|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C700-C701,C709|Meninges|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C700-C701,C709|Meninges|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C700-C701,C709|Meninges|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C700-C701,C709|Meninges|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C700-C701,C709|Meninges|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C700-C701,C709|Meninges|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C700-C701,C709|Meninges|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C700-C701,C709|Meninges|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C700-C701,C709|Meninges|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C700-C701,C709|Meninges|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C700-C701,C709|Meninges|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C700-C701,C709|Meninges|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C700-C701,C709|Meninges|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C700-C701,C709|Meninges|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C700-C701,C709|Meninges|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9812/3|null
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9813/3|null
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9814/3|null
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9817/3|null
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9818/3|null
C700-C701,C709|Meninges|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C700-C701,C709|Meninges|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C700-C701,C709|Meninges|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C700-C701,C709|Meninges|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C700-C701,C709|Meninges|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C700-C701,C709|Meninges|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C700-C701,C709|Meninges|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C700-C701,C709|Meninges|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C710-C714, C717-C719, C720-C725|CranialNerve|868|Paraganglioma|8680/1|Paraganglioma
C710-C714, C717-C719, C720-C725|CranialNerve|872|Melanoma|8720/3|Melanoma
C710-C714, C717-C719, C720-C725|CranialNerve|880|Sarcoma|8800/0|BenignSoftTissueNeoplasm
C710-C714, C717-C719, C720-C725|CranialNerve|880|Sarcoma|8800/3|Sarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|880|Sarcoma|8801/3|SpindleCellSarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C710-C714, C717-C719, C720-C725|CranialNerve|881|FibromatousNeoplasm|8815/1|null
C710-C714, C717-C719, C720-C725|CranialNerve|881|FibromatousNeoplasm|8815/3|MalignantHemangiopericytoma
C710-C714, C717-C719, C720-C725|CranialNerve|885|Liposarcoma|8850/0|Lipoma
C710-C714, C717-C719, C720-C725|CranialNerve|885|Liposarcoma|8851/0|Fibrolipoma
C710-C714, C717-C719, C720-C725|CranialNerve|885|Liposarcoma|8851/3|WellDifferentiatedLiposarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|906|GermCellTumor|9060/3|Dysgerminoma
C710-C714, C717-C719, C720-C725|CranialNerve|906|GermCellTumor|9064/3|Germinoma
C710-C714, C717-C719, C720-C725|CranialNerve|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C710-C714, C717-C719, C720-C725|CranialNerve|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C710-C714, C717-C719, C720-C725|CranialNerve|908|Teratoma|9080/0|MatureTeratoma
C710-C714, C717-C719, C720-C725|CranialNerve|908|Teratoma|9080/1|Teratoma
C710-C714, C717-C719, C720-C725|CranialNerve|908|Teratoma|9080/3|ImmatureTeratoma
C710-C714, C717-C719, C720-C725|CranialNerve|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C710-C714, C717-C719, C720-C725|CranialNerve|908|Teratoma|9085/3|MixedGermCellTumor
C710-C714, C717-C719, C720-C725|CranialNerve|910|Choriocarcinoma|9100/3|Choriocarcinoma
C710-C714, C717-C719, C720-C725|CranialNerve|912|NeoplasmsVascularTissue|9120/0|Hemangioma
C710-C714, C717-C719, C720-C725|CranialNerve|912|NeoplasmsVascularTissue|9121/0|HemangiomaCavernous
C710-C714, C717-C719, C720-C725|CranialNerve|912|NeoplasmsVascularTissue|9122/0|VenousHemangioma
C710-C714, C717-C719, C720-C725|CranialNerve|913|Hemangioendothelioma|9131/0|CapillaryHemangioma
C710-C714, C717-C719, C720-C725|CranialNerve|915|Hemangiopericytoma|9150/1|Hemangiopericytoma
C710-C714, C717-C719, C720-C725|CranialNerve|916|Hemangioblastoma|9161/1|Hemangioblastoma
C710-C714, C717-C719, C720-C725|CranialNerve|937|Chordoma|9370/3|Chordoma
C710-C714, C717-C719, C720-C725|CranialNerve|937|Chordoma|9371/3|ChondroidChordoma
C710-C714, C717-C719, C720-C725|CranialNerve|937|Chordoma|9372/3|DedifferentiatedChordoma
C710-C714, C717-C719, C720-C725|CranialNerve|938|Glioma|9380/1|Glioma
C710-C714, C717-C719, C720-C725|CranialNerve|938|Glioma|9380/3|MalignantGlioma
C710-C714, C717-C719, C720-C725|CranialNerve|938|Glioma|9381/3|GliomatosisCerebri
C710-C714, C717-C719, C720-C725|CranialNerve|938|Glioma|9382/3|MixedGlioma
C710-C714, C717-C719, C720-C725|CranialNerve|938|Glioma|9383/1|SubependymalGlioma
C710-C714, C717-C719, C720-C725|CranialNerve|938|Glioma|9384/1|Astrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|938|Glioma|9385/3|Glioma
C710-C714, C717-C719, C720-C725|CranialNerve|939|Ependymoma|9391/3|Ependymoma
C710-C714, C717-C719, C720-C725|CranialNerve|939|Ependymoma|9392/3|AnaplasticEpendymoma
C710-C714, C717-C719, C720-C725|CranialNerve|939|Ependymoma|9393/3|PapillaryEpendymoma
C710-C714, C717-C719, C720-C725|CranialNerve|939|Ependymoma|9394/1|MyxopapillaryEpendymoma
C710-C714, C717-C719, C720-C725|CranialNerve|939|Ependymoma|9396/3|EpendymomaRELAFusionPositive
C710-C714, C717-C719, C720-C725|CranialNerve|940|Astrocytoma|9400/3|Astrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|940|Astrocytoma|9401/3|AnaplasticAstrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|941|ProtoplasmicAstrocytoma|9410/3|ProtoplasmicAstrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|941|ProtoplasmicAstrocytoma|9411/3|GemistocyticAstrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|941|ProtoplasmicAstrocytoma|9412/1|DesmoplasticInfantileAstrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|941|ProtoplasmicAstrocytoma|9413/0|DysembryoplasticNeuroepithelialTumor
C710-C714, C717-C719, C720-C725|CranialNerve|942|FibrillaryAstrocytoma|9420/3|FibrillaryAstrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|942|FibrillaryAstrocytoma|9421/1|PilocyticAstrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|942|FibrillaryAstrocytoma|9421/3|PilocyticAstrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|942|FibrillaryAstrocytoma|9423/3|PolarSpongioblastoma
C710-C714, C717-C719, C720-C725|CranialNerve|942|FibrillaryAstrocytoma|9424/3|PleomorphicXanthoastrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|942|FibrillaryAstrocytoma|9425/3|PilomyxoidAstrocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|943|Astroblastoma|9430/3|Astroblastoma
C710-C714, C717-C719, C720-C725|CranialNerve|943|Astroblastoma|9431/1|AngiocentricGlioma
C710-C714, C717-C719, C720-C725|CranialNerve|944|Glioblastoma|9440/1|BrainNeoplasm
C710-C714, C717-C719, C720-C725|CranialNerve|944|Glioblastoma|9440/3|Glioblastoma
C710-C714, C717-C719, C720-C725|CranialNerve|944|Glioblastoma|9441/3|GiantCellGlioblastoma
C710-C714, C717-C719, C720-C725|CranialNerve|944|Glioblastoma|9442/1|Gliofibroma
C710-C714, C717-C719, C720-C725|CranialNerve|944|Glioblastoma|9442/3|Gliosarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|944|Glioblastoma|9444/1|ChordoidGliomaOfTheThirdVentricle
C710-C714, C717-C719, C720-C725|CranialNerve|944|Glioblastoma|9445/3|GlioblastomaIDHMutant
C710-C714, C717-C719, C720-C725|CranialNerve|945|AdultOligodendroglioma|9450/3|AdultOligodendroglioma
C710-C714, C717-C719, C720-C725|CranialNerve|945|AdultOligodendroglioma|9451/3|AnaplasticOligodendroglioma
C710-C714, C717-C719, C720-C725|CranialNerve|946|Oligodendroblastoma|9460/3|Oligodendroblastoma
C710-C714, C717-C719, C720-C725|CranialNerve|947|Medulloblastoma|9473/3|PrimitiveNeuroectodermalTumor
C710-C714, C717-C719, C720-C725|CranialNerve|947|Medulloblastoma|9475/3|MedulloblastomaWNTActivated
C710-C714, C717-C719, C720-C725|CranialNerve|947|Medulloblastoma|9476/3|MedulloblastomaSHHActivated
C710-C714, C717-C719, C720-C725|CranialNerve|947|Medulloblastoma|9477/3|MedulloblastomaNonWNTNonSHH
C710-C714, C717-C719, C720-C725|CranialNerve|947|Medulloblastoma|9478/3|EmbryonalNeoplasm
C710-C714, C717-C719, C720-C725|CranialNerve|949|Ganglioneuroblastoma|9490/0|Ganglioneuroma
C710-C714, C717-C719, C720-C725|CranialNerve|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C710-C714, C717-C719, C720-C725|CranialNerve|949|Ganglioneuroblastoma|9492/0|Gangliocytoma
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9500/3|Neuroblastoma
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9501/3|Medulloepithelioma
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9503/3|Neuroepithelioma
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9505/0|NeuronalChoristoma
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9505/1|Ganglioglioma
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9508/3|AtypicalTeratoidRhabdoidTumorCL372028
C710-C714, C717-C719, C720-C725|CranialNerve|950|Neuroblastoma|9509/1|PapillaryGlioneuronalTumor
C710-C714, C717-C719, C720-C725|CranialNerve|954|MalignantPeripheralNerveSheathTumor|9540/0|Neurofibroma
C710-C714, C717-C719, C720-C725|CranialNerve|954|MalignantPeripheralNerveSheathTumor|9540/1|Neurofibromatosis
C710-C714, C717-C719, C720-C725|CranialNerve|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C710-C714, C717-C719, C720-C725|CranialNerve|954|MalignantPeripheralNerveSheathTumor|9541/0|MelanoticNeurofibroma
C710-C714, C717-C719, C720-C725|CranialNerve|955|PlexiformNeurofibroma|9550/0|PlexiformNeurofibroma
C710-C714, C717-C719, C720-C725|CranialNerve|956|Schwannoma|9560/0|Schwannoma
C710-C714, C717-C719, C720-C725|CranialNerve|956|Schwannoma|9560/1|MelanoticSchwannoma
C710-C714, C717-C719, C720-C725|CranialNerve|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C710-C714, C717-C719, C720-C725|CranialNerve|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C710-C714, C717-C719, C720-C725|CranialNerve|956|Schwannoma|9562/0|Neurothekeoma
C710-C714, C717-C719, C720-C725|CranialNerve|957|Perineurioma|9570/0|Neuroma
C710-C714, C717-C719, C720-C725|CranialNerve|957|Perineurioma|9571/0|Perineurioma
C710-C714, C717-C719, C720-C725|CranialNerve|957|Perineurioma|9571/3|MalignantPerineurioma
C710-C714, C717-C719, C720-C725|CranialNerve|959|Lymphoma|9590/3|Lymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|959|Lymphoma|9596/3|CompositeLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|967|BCellLymphomas|9673/3|MantleCellLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|969|FollicularAdenoma|9690/3|LymphomaFollicular
C710-C714, C717-C719, C720-C725|CranialNerve|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C710-C714, C717-C719, C720-C725|CranialNerve|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C710-C714, C717-C719, C720-C725|CranialNerve|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|970|TCellLymphoma|9701/3|SezarySyndrome
C710-C714, C717-C719, C720-C725|CranialNerve|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C710-C714, C717-C719, C720-C725|CranialNerve|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C710-C714, C717-C719, C720-C725|CranialNerve|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C710-C714, C717-C719, C720-C725|CranialNerve|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C710-C714, C717-C719, C720-C725|CranialNerve|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C710-C714, C717-C719, C720-C725|CranialNerve|973|Plasmacytoma|9731/3|Plasmacytoma
C710-C714, C717-C719, C720-C725|CranialNerve|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C710-C714, C717-C719, C720-C725|CranialNerve|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C710-C714, C717-C719, C720-C725|CranialNerve|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C710-C714, C717-C719, C720-C725|CranialNerve|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C710-C714, C717-C719, C720-C725|CranialNerve|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C710-C714, C717-C719, C720-C725|CranialNerve|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C710-C714, C717-C719, C720-C725|CranialNerve|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C710-C714, C717-C719, C720-C725|CranialNerve|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9812/3|null
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9813/3|null
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9814/3|null
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9817/3|null
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9818/3|null
C710-C714, C717-C719, C720-C725|CranialNerve|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C710-C714, C717-C719, C720-C725|CranialNerve|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C710-C714, C717-C719, C720-C725|CranialNerve|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C710-C714, C717-C719, C720-C725|CranialNerve|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C710-C714, C717-C719, C720-C725|CranialNerve|993|MyeloidSarcoma|9930/3|MyeloidSarcoma
C710-C714, C717-C719, C720-C725|CranialNerve|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C710-C714, C717-C719, C720-C725|CranialNerve|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C710-C714, C717-C719, C720-C725|CranialNerve|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C710-C714, C717-C719, C720-C725|CranialNerve|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C715|BrainVentricle|908|Teratoma|9085/3|MixedGermCellTumor
C715|BrainVentricle|937|Chordoma|9370/3|Chordoma
C715|BrainVentricle|937|Chordoma|9371/3|ChondroidChordoma
C715|BrainVentricle|937|Chordoma|9372/3|DedifferentiatedChordoma
C715|BrainVentricle|938|Glioma|9380/3|MalignantGlioma
C715|BrainVentricle|938|Glioma|9381/3|GliomatosisCerebri
C715|BrainVentricle|938|Glioma|9382/3|MixedGlioma
C715|BrainVentricle|938|Glioma|9383/1|SubependymalGlioma
C715|BrainVentricle|938|Glioma|9384/1|Astrocytoma
C715|BrainVentricle|938|Glioma|9385/3|Glioma
C715|BrainVentricle|939|Ependymoma|9390/0|ChoroidPlexusPapilloma
C715|BrainVentricle|939|Ependymoma|9390/1|AtypicalChoroidPlexusPapilloma
C715|BrainVentricle|939|Ependymoma|9390/3|ChoroidPlexusCarcinoma
C715|BrainVentricle|939|Ependymoma|9391/3|Ependymoma
C715|BrainVentricle|939|Ependymoma|9392/3|AnaplasticEpendymoma
C715|BrainVentricle|939|Ependymoma|9393/3|PapillaryEpendymoma
C715|BrainVentricle|939|Ependymoma|9396/3|EpendymomaRELAFusionPositive
C715|BrainVentricle|940|Astrocytoma|9400/3|Astrocytoma
C715|BrainVentricle|940|Astrocytoma|9401/3|AnaplasticAstrocytoma
C715|BrainVentricle|941|ProtoplasmicAstrocytoma|9410/3|ProtoplasmicAstrocytoma
C715|BrainVentricle|941|ProtoplasmicAstrocytoma|9411/3|GemistocyticAstrocytoma
C715|BrainVentricle|942|FibrillaryAstrocytoma|9420/3|FibrillaryAstrocytoma
C715|BrainVentricle|942|FibrillaryAstrocytoma|9421/1|PilocyticAstrocytoma
C715|BrainVentricle|942|FibrillaryAstrocytoma|9421/3|PilocyticAstrocytoma
C715|BrainVentricle|942|FibrillaryAstrocytoma|9423/3|PolarSpongioblastoma
C715|BrainVentricle|942|FibrillaryAstrocytoma|9424/3|PleomorphicXanthoastrocytoma
C715|BrainVentricle|942|FibrillaryAstrocytoma|9425/3|PilomyxoidAstrocytoma
C715|BrainVentricle|943|Astroblastoma|9430/3|Astroblastoma
C715|BrainVentricle|943|Astroblastoma|9431/1|AngiocentricGlioma
C715|BrainVentricle|944|Glioblastoma|9440/3|Glioblastoma
C715|BrainVentricle|944|Glioblastoma|9441/3|GiantCellGlioblastoma
C715|BrainVentricle|944|Glioblastoma|9442/3|Gliosarcoma
C715|BrainVentricle|944|Glioblastoma|9444/1|ChordoidGliomaOfTheThirdVentricle
C715|BrainVentricle|944|Glioblastoma|9445/3|GlioblastomaIDHMutant
C715|BrainVentricle|945|AdultOligodendroglioma|9450/3|AdultOligodendroglioma
C715|BrainVentricle|945|AdultOligodendroglioma|9451/3|AnaplasticOligodendroglioma
C715|BrainVentricle|947|Medulloblastoma|9473/3|PrimitiveNeuroectodermalTumor
C715|BrainVentricle|947|Medulloblastoma|9475/3|MedulloblastomaWNTActivated
C715|BrainVentricle|947|Medulloblastoma|9476/3|MedulloblastomaSHHActivated
C715|BrainVentricle|947|Medulloblastoma|9477/3|MedulloblastomaNonWNTNonSHH
C715|BrainVentricle|947|Medulloblastoma|9478/3|EmbryonalNeoplasm
C715|BrainVentricle|949|Ganglioneuroblastoma|9490/0|Ganglioneuroma
C715|BrainVentricle|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C715|BrainVentricle|949|Ganglioneuroblastoma|9492/0|Gangliocytoma
C715|BrainVentricle|950|Neuroblastoma|9500/3|Neuroblastoma
C715|BrainVentricle|950|Neuroblastoma|9501/3|Medulloepithelioma
C715|BrainVentricle|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C715|BrainVentricle|950|Neuroblastoma|9503/3|Neuroepithelioma
C715|BrainVentricle|950|Neuroblastoma|9505/1|Ganglioglioma
C715|BrainVentricle|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C715|BrainVentricle|950|Neuroblastoma|9506/1|Neurocytoma
C715|BrainVentricle|950|Neuroblastoma|9508/3|AtypicalTeratoidRhabdoidTumorCL372028
C715|BrainVentricle|950|Neuroblastoma|9509/1|PapillaryGlioneuronalTumor
C715|BrainVentricle|959|Lymphoma|9590/3|Lymphoma
C715|BrainVentricle|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C715|BrainVentricle|959|Lymphoma|9596/3|CompositeLymphoma
C715|BrainVentricle|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C715|BrainVentricle|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C715|BrainVentricle|967|BCellLymphomas|9673/3|MantleCellLymphoma
C715|BrainVentricle|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C715|BrainVentricle|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C715|BrainVentricle|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C715|BrainVentricle|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C715|BrainVentricle|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C715|BrainVentricle|969|FollicularAdenoma|9690/3|LymphomaFollicular
C715|BrainVentricle|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C715|BrainVentricle|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C715|BrainVentricle|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C715|BrainVentricle|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C715|BrainVentricle|970|TCellLymphoma|9701/3|SezarySyndrome
C715|BrainVentricle|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C715|BrainVentricle|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C715|BrainVentricle|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C715|BrainVentricle|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C715|BrainVentricle|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C715|BrainVentricle|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C715|BrainVentricle|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C715|BrainVentricle|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C715|BrainVentricle|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C715|BrainVentricle|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C715|BrainVentricle|973|Plasmacytoma|9731/3|Plasmacytoma
C715|BrainVentricle|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C715|BrainVentricle|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C715|BrainVentricle|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C715|BrainVentricle|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C715|BrainVentricle|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C715|BrainVentricle|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C715|BrainVentricle|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C715|BrainVentricle|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C715|BrainVentricle|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C715|BrainVentricle|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C715|BrainVentricle|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C715|BrainVentricle|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C715|BrainVentricle|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C715|BrainVentricle|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9812/3|null
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9813/3|null
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9814/3|null
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9817/3|null
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9818/3|null
C715|BrainVentricle|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C715|BrainVentricle|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C715|BrainVentricle|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C715|BrainVentricle|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C715|BrainVentricle|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C715|BrainVentricle|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C715|BrainVentricle|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C715|BrainVentricle|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C716|Cerebellum|880|Sarcoma|8800/0|BenignSoftTissueNeoplasm
C716|Cerebellum|880|Sarcoma|8800/3|Sarcoma
C716|Cerebellum|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C716|Cerebellum|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C716|Cerebellum|881|FibromatousNeoplasm|8810/3|Fibrosarcoma
C716|Cerebellum|881|FibromatousNeoplasm|8815/0|SolitaryFibrousTumor
C716|Cerebellum|882|Sarcoma|8825/3|LowGradeMyofibroblasticSarcoma
C716|Cerebellum|885|Liposarcoma|8850/0|Lipoma
C716|Cerebellum|908|Teratoma|9080/0|MatureTeratoma
C716|Cerebellum|908|Teratoma|9080/1|Teratoma
C716|Cerebellum|908|Teratoma|9080/3|ImmatureTeratoma
C716|Cerebellum|908|Teratoma|9084/0|DermoidCyst
C716|Cerebellum|912|NeoplasmsVascularTissue|9120/0|Hemangioma
C716|Cerebellum|913|Hemangioendothelioma|9131/0|CapillaryHemangioma
C716|Cerebellum|915|Hemangiopericytoma|9150/1|Hemangiopericytoma
C716|Cerebellum|916|Hemangioblastoma|9161/1|Hemangioblastoma
C716|Cerebellum|937|Chordoma|9370/3|Chordoma
C716|Cerebellum|937|Chordoma|9371/3|ChondroidChordoma
C716|Cerebellum|937|Chordoma|9372/3|DedifferentiatedChordoma
C716|Cerebellum|938|Glioma|9380/1|Glioma
C716|Cerebellum|938|Glioma|9380/3|MalignantGlioma
C716|Cerebellum|938|Glioma|9381/3|GliomatosisCerebri
C716|Cerebellum|938|Glioma|9382/3|MixedGlioma
C716|Cerebellum|938|Glioma|9383/1|SubependymalGlioma
C716|Cerebellum|938|Glioma|9385/3|Glioma
C716|Cerebellum|939|Ependymoma|9391/3|Ependymoma
C716|Cerebellum|939|Ependymoma|9392/3|AnaplasticEpendymoma
C716|Cerebellum|939|Ependymoma|9393/3|PapillaryEpendymoma
C716|Cerebellum|939|Ependymoma|9396/3|EpendymomaRELAFusionPositive
C716|Cerebellum|940|Astrocytoma|9400/3|Astrocytoma
C716|Cerebellum|940|Astrocytoma|9401/3|AnaplasticAstrocytoma
C716|Cerebellum|941|ProtoplasmicAstrocytoma|9410/3|ProtoplasmicAstrocytoma
C716|Cerebellum|941|ProtoplasmicAstrocytoma|9411/3|GemistocyticAstrocytoma
C716|Cerebellum|942|FibrillaryAstrocytoma|9420/3|FibrillaryAstrocytoma
C716|Cerebellum|942|FibrillaryAstrocytoma|9421/1|PilocyticAstrocytoma
C716|Cerebellum|942|FibrillaryAstrocytoma|9421/3|PilocyticAstrocytoma
C716|Cerebellum|942|FibrillaryAstrocytoma|9424/3|PleomorphicXanthoastrocytoma
C716|Cerebellum|942|FibrillaryAstrocytoma|9425/3|PilomyxoidAstrocytoma
C716|Cerebellum|943|Astroblastoma|9430/3|Astroblastoma
C716|Cerebellum|943|Astroblastoma|9431/1|AngiocentricGlioma
C716|Cerebellum|944|Glioblastoma|9440/3|Glioblastoma
C716|Cerebellum|944|Glioblastoma|9441/3|GiantCellGlioblastoma
C716|Cerebellum|944|Glioblastoma|9442/3|Gliosarcoma
C716|Cerebellum|944|Glioblastoma|9445/3|GlioblastomaIDHMutant
C716|Cerebellum|945|AdultOligodendroglioma|9450/3|AdultOligodendroglioma
C716|Cerebellum|945|AdultOligodendroglioma|9451/3|AnaplasticOligodendroglioma
C716|Cerebellum|947|Medulloblastoma|9470/3|Medulloblastoma
C716|Cerebellum|947|Medulloblastoma|9471/3|DesmoplasticNodularMedulloblastoma
C716|Cerebellum|947|Medulloblastoma|9472/3|Medullomyoblastoma
C716|Cerebellum|947|Medulloblastoma|9473/3|PrimitiveNeuroectodermalTumor
C716|Cerebellum|947|Medulloblastoma|9474/3|LargeCellMedulloblastoma
C716|Cerebellum|947|Medulloblastoma|9475/3|MedulloblastomaWNTActivated
C716|Cerebellum|947|Medulloblastoma|9476/3|MedulloblastomaSHHActivated
C716|Cerebellum|947|Medulloblastoma|9477/3|MedulloblastomaNonWNTNonSHH
C716|Cerebellum|947|Medulloblastoma|9478/3|EmbryonalNeoplasm
C716|Cerebellum|948|CerebellarSarcoma|9480/3|CerebellarSarcoma
C716|Cerebellum|949|Ganglioneuroblastoma|9490/0|Ganglioneuroma
C716|Cerebellum|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C716|Cerebellum|949|Ganglioneuroblastoma|9492/0|Gangliocytoma
C716|Cerebellum|949|Ganglioneuroblastoma|9493/0|LhermitteDuclosDisease
C716|Cerebellum|950|Neuroblastoma|9500/3|Neuroblastoma
C716|Cerebellum|950|Neuroblastoma|9501/3|Medulloepithelioma
C716|Cerebellum|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C716|Cerebellum|950|Neuroblastoma|9503/3|Neuroepithelioma
C716|Cerebellum|950|Neuroblastoma|9505/1|Ganglioglioma
C716|Cerebellum|950|Neuroblastoma|9506/1|Neurocytoma
C716|Cerebellum|950|Neuroblastoma|9508/3|AtypicalTeratoidRhabdoidTumorCL372028
C716|Cerebellum|950|Neuroblastoma|9509/1|PapillaryGlioneuronalTumor
C716|Cerebellum|959|Lymphoma|9590/3|Lymphoma
C716|Cerebellum|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C716|Cerebellum|959|Lymphoma|9596/3|CompositeLymphoma
C716|Cerebellum|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C716|Cerebellum|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C716|Cerebellum|967|BCellLymphomas|9673/3|MantleCellLymphoma
C716|Cerebellum|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C716|Cerebellum|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C716|Cerebellum|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C716|Cerebellum|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C716|Cerebellum|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C716|Cerebellum|969|FollicularAdenoma|9690/3|LymphomaFollicular
C716|Cerebellum|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C716|Cerebellum|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C716|Cerebellum|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C716|Cerebellum|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C716|Cerebellum|970|TCellLymphoma|9701/3|SezarySyndrome
C716|Cerebellum|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C716|Cerebellum|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C716|Cerebellum|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C716|Cerebellum|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C716|Cerebellum|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C716|Cerebellum|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C716|Cerebellum|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C716|Cerebellum|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C716|Cerebellum|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C716|Cerebellum|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C716|Cerebellum|973|Plasmacytoma|9731/3|Plasmacytoma
C716|Cerebellum|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C716|Cerebellum|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C716|Cerebellum|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C716|Cerebellum|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C716|Cerebellum|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C716|Cerebellum|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C716|Cerebellum|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C716|Cerebellum|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C716|Cerebellum|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C716|Cerebellum|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C716|Cerebellum|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C716|Cerebellum|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C716|Cerebellum|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C716|Cerebellum|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9812/3|null
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9813/3|null
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9814/3|null
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9817/3|null
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9818/3|null
C716|Cerebellum|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C716|Cerebellum|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C716|Cerebellum|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C716|Cerebellum|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C716|Cerebellum|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C716|Cerebellum|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C716|Cerebellum|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C716|Cerebellum|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C728-C729|CentralNervousSystem|880|Sarcoma|8800/0|BenignSoftTissueNeoplasm
C728-C729|CentralNervousSystem|880|Sarcoma|8800/3|Sarcoma
C728-C729|CentralNervousSystem|880|Sarcoma|8801/3|SpindleCellSarcoma
C728-C729|CentralNervousSystem|880|Sarcoma|8802/3|GiantCellSarcoma
C728-C729|CentralNervousSystem|880|Sarcoma|8803/3|SmallCellSarcoma
C728-C729|CentralNervousSystem|880|Sarcoma|8804/3|SarcomaEpithelioid
C728-C729|CentralNervousSystem|880|Sarcoma|8805/3|UndifferentiatedSarcoma
C728-C729|CentralNervousSystem|880|Sarcoma|8806/3|DesmoplasticSmallRoundCellTumor
C728-C729|CentralNervousSystem|885|Liposarcoma|8850/0|Lipoma
C728-C729|CentralNervousSystem|885|Liposarcoma|8850/1|AtypicalLipoma
C728-C729|CentralNervousSystem|885|Liposarcoma|8850/3|Liposarcoma
C728-C729|CentralNervousSystem|886|Angiolipoma|8861/0|Angiolipoma
C728-C729|CentralNervousSystem|889|MyomatousNeoplasm|8890/0|FibroidTumor
C728-C729|CentralNervousSystem|889|MyomatousNeoplasm|8890/1|Leiomyomatosis
C728-C729|CentralNervousSystem|889|MyomatousNeoplasm|8890/3|Leiomyosarcoma
C728-C729|CentralNervousSystem|889|MyomatousNeoplasm|8897/1|SmoothMuscleNeoplasm
C728-C729|CentralNervousSystem|890|Rhabdomyosarcoma|8900/0|Rhabdomyoma
C728-C729|CentralNervousSystem|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C728-C729|CentralNervousSystem|891|EmbryonalRhabdomyosarcoma|8910/3|EmbryonalRhabdomyosarcoma
C728-C729|CentralNervousSystem|892|AlveolarRhabdomyosarcoma|8920/3|AlveolarRhabdomyosarcoma
C728-C729|CentralNervousSystem|906|GermCellTumor|9064/3|Germinoma
C728-C729|CentralNervousSystem|908|Teratoma|9080/1|Teratoma
C728-C729|CentralNervousSystem|908|Teratoma|9080/3|ImmatureTeratoma
C728-C729|CentralNervousSystem|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C728-C729|CentralNervousSystem|908|Teratoma|9084/0|DermoidCyst
C728-C729|CentralNervousSystem|908|Teratoma|9084/3|Teratoma
C728-C729|CentralNervousSystem|912|NeoplasmsVascularTissue|9120/0|Hemangioma
C728-C729|CentralNervousSystem|912|NeoplasmsVascularTissue|9120/3|Hemangiosarcoma
C728-C729|CentralNervousSystem|912|NeoplasmsVascularTissue|9121/0|HemangiomaCavernous
C728-C729|CentralNervousSystem|913|Hemangioendothelioma|9130/0|BenignHemangioendothelioma
C728-C729|CentralNervousSystem|913|Hemangioendothelioma|9130/1|Hemangioendothelioma
C728-C729|CentralNervousSystem|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C728-C729|CentralNervousSystem|914|KaposiSarcoma|9140/3|KaposiSarcoma
C728-C729|CentralNervousSystem|915|Hemangiopericytoma|9150/0|BenignHemangiopericytoma
C728-C729|CentralNervousSystem|915|Hemangiopericytoma|9150/1|Hemangiopericytoma
C728-C729|CentralNervousSystem|915|Hemangiopericytoma|9150/3|MalignantHemangiopericytoma
C728-C729|CentralNervousSystem|916|Hemangioblastoma|9161/1|Hemangioblastoma
C728-C729|CentralNervousSystem|926|EwingSarcoma|9260/3|EwingSarcoma
C728-C729|CentralNervousSystem|937|Chordoma|9370/3|Chordoma
C728-C729|CentralNervousSystem|937|Chordoma|9371/3|ChondroidChordoma
C728-C729|CentralNervousSystem|937|Chordoma|9372/3|DedifferentiatedChordoma
C728-C729|CentralNervousSystem|950|Neuroblastoma|9500/3|Neuroblastoma
C728-C729|CentralNervousSystem|950|Neuroblastoma|9501/3|Medulloepithelioma
C728-C729|CentralNervousSystem|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C728-C729|CentralNervousSystem|950|Neuroblastoma|9503/3|Neuroepithelioma
C728-C729|CentralNervousSystem|950|Neuroblastoma|9508/3|AtypicalTeratoidRhabdoidTumorCL372028
C728-C729|CentralNervousSystem|954|MalignantPeripheralNerveSheathTumor|9540/0|Neurofibroma
C728-C729|CentralNervousSystem|954|MalignantPeripheralNerveSheathTumor|9540/1|Neurofibromatosis
C728-C729|CentralNervousSystem|954|MalignantPeripheralNerveSheathTumor|9540/3|MalignantPeripheralNerveSheathTumor
C728-C729|CentralNervousSystem|954|MalignantPeripheralNerveSheathTumor|9541/0|MelanoticNeurofibroma
C728-C729|CentralNervousSystem|955|PlexiformNeurofibroma|9550/0|PlexiformNeurofibroma
C728-C729|CentralNervousSystem|956|Schwannoma|9560/0|Schwannoma
C728-C729|CentralNervousSystem|956|Schwannoma|9560/3|MalignantPeripheralNerveSheathTumor
C728-C729|CentralNervousSystem|956|Schwannoma|9561/3|MalignantPeripheralNerveSheathTumor
C728-C729|CentralNervousSystem|956|Schwannoma|9562/0|Neurothekeoma
C728-C729|CentralNervousSystem|957|Perineurioma|9570/0|Neuroma
C728-C729|CentralNervousSystem|957|Perineurioma|9571/0|Perineurioma
C728-C729|CentralNervousSystem|957|Perineurioma|9571/3|MalignantPerineurioma
C728-C729|CentralNervousSystem|959|Lymphoma|9590/3|Lymphoma
C728-C729|CentralNervousSystem|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C728-C729|CentralNervousSystem|959|Lymphoma|9596/3|CompositeLymphoma
C728-C729|CentralNervousSystem|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C728-C729|CentralNervousSystem|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C728-C729|CentralNervousSystem|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C728-C729|CentralNervousSystem|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C728-C729|CentralNervousSystem|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C728-C729|CentralNervousSystem|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C728-C729|CentralNervousSystem|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C728-C729|CentralNervousSystem|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C728-C729|CentralNervousSystem|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C728-C729|CentralNervousSystem|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C728-C729|CentralNervousSystem|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C728-C729|CentralNervousSystem|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C728-C729|CentralNervousSystem|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C728-C729|CentralNervousSystem|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C728-C729|CentralNervousSystem|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C728-C729|CentralNervousSystem|967|BCellLymphomas|9673/3|MantleCellLymphoma
C728-C729|CentralNervousSystem|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C728-C729|CentralNervousSystem|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C728-C729|CentralNervousSystem|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C728-C729|CentralNervousSystem|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C728-C729|CentralNervousSystem|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C728-C729|CentralNervousSystem|969|FollicularAdenoma|9690/3|LymphomaFollicular
C728-C729|CentralNervousSystem|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C728-C729|CentralNervousSystem|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C728-C729|CentralNervousSystem|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C728-C729|CentralNervousSystem|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C728-C729|CentralNervousSystem|970|TCellLymphoma|9701/3|SezarySyndrome
C728-C729|CentralNervousSystem|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C728-C729|CentralNervousSystem|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C728-C729|CentralNervousSystem|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C728-C729|CentralNervousSystem|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C728-C729|CentralNervousSystem|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C728-C729|CentralNervousSystem|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C728-C729|CentralNervousSystem|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C728-C729|CentralNervousSystem|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C728-C729|CentralNervousSystem|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C728-C729|CentralNervousSystem|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C728-C729|CentralNervousSystem|973|Plasmacytoma|9731/3|Plasmacytoma
C728-C729|CentralNervousSystem|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C728-C729|CentralNervousSystem|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C728-C729|CentralNervousSystem|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C728-C729|CentralNervousSystem|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C728-C729|CentralNervousSystem|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C728-C729|CentralNervousSystem|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C728-C729|CentralNervousSystem|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C728-C729|CentralNervousSystem|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C728-C729|CentralNervousSystem|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C728-C729|CentralNervousSystem|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C728-C729|CentralNervousSystem|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C728-C729|CentralNervousSystem|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C728-C729|CentralNervousSystem|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C728-C729|CentralNervousSystem|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C728-C729|CentralNervousSystem|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C728-C729|CentralNervousSystem|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9812/3|null
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9813/3|null
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9814/3|null
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9817/3|null
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9818/3|null
C728-C729|CentralNervousSystem|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C728-C729|CentralNervousSystem|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C728-C729|CentralNervousSystem|982|LymphoidLeukemia|9827/3|AdultTcellLeukemia
C728-C729|CentralNervousSystem|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C728-C729|CentralNervousSystem|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C728-C729|CentralNervousSystem|986|MyeloidLeukemia|9861/3|AcuteMyeloidLeukemia
C728-C729|CentralNervousSystem|993|MyeloidSarcoma|9930/3|MyeloidSarcoma
C728-C729|CentralNervousSystem|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C728-C729|CentralNervousSystem|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C728-C729|CentralNervousSystem|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C728-C729|CentralNervousSystem|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C739|ThyroidGland|801|Carcinoma|8010/2|InSituCancer
C739|ThyroidGland|801|Carcinoma|8010/3|CarcinomaNOSDNE
C739|ThyroidGland|801|Carcinoma|8011/3|MalignantEpithelioma
C739|ThyroidGland|801|Carcinoma|8012/3|LargeCellCarcinoma
C739|ThyroidGland|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C739|ThyroidGland|801|Carcinoma|8014/3|LargeCellCarcinoma
C739|ThyroidGland|801|Carcinoma|8015/3|GlassyCellCarcinoma
C739|ThyroidGland|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C739|ThyroidGland|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C739|ThyroidGland|802|Carcinoma|8022/3|PleomorphicCarcinoma
C739|ThyroidGland|803|SarcomatoidCarcinoma|8030/3|GiantCellAndSpindleCellCarcinoma
C739|ThyroidGland|803|SarcomatoidCarcinoma|8031/3|GiantCellCarcinoma
C739|ThyroidGland|803|SarcomatoidCarcinoma|8032/3|SarcomatoidCarcinoma
C739|ThyroidGland|803|SarcomatoidCarcinoma|8033/3|SarcomatoidCarcinoma
C739|ThyroidGland|803|SarcomatoidCarcinoma|8034/3|PolygonalCellCarcinoma
C739|ThyroidGland|803|SarcomatoidCarcinoma|8035/3|NeoplasticOsteoclastLikeGiantCell
C739|ThyroidGland|804|SmallCellCarcinoma|8041/3|SmallCellCarcinoma
C739|ThyroidGland|804|SmallCellCarcinoma|8041/6|MetastaticSmallCellCarcinoma
C739|ThyroidGland|804|SmallCellCarcinoma|8043/3|SmallCellCarcinomaFusiformCell
C739|ThyroidGland|805|PapillaryCarcinoma|8050/2|PapillaryCarcinomaInSitu
C739|ThyroidGland|805|PapillaryCarcinoma|8050/3|PapillaryCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8070/2|Stage0SquamousCellCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8070/3|SquamousCellCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8071/3|KeratinizingMalignantSquamousCell
C739|ThyroidGland|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8072/3|NonkeratinisingSquamousCellCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8074/3|SarcomatoidCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8075/3|PseudoglandularSquamousCellCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8076/2|Stage0SquamousCellCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8076/3|MicroinvasiveSquamousCellCarcinoma
C739|ThyroidGland|807|SquamousCellCarcinoma|8078/3|MicroinvasiveSquamousCellCarcinoma
C739|ThyroidGland|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C739|ThyroidGland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C739|ThyroidGland|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C739|ThyroidGland|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C739|ThyroidGland|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C739|ThyroidGland|819|TrabecularAdenocarcinoma|8190/3|TrabecularAdenocarcinoma
C739|ThyroidGland|823|SolidCarcinoma|8230/2|InSituCancer
C739|ThyroidGland|823|SolidCarcinoma|8230/3|SolidCarcinoma
C739|ThyroidGland|823|SolidCarcinoma|8231/3|CarcinomaSimplex
C739|ThyroidGland|825|BronchioloalveolarAdenocarcinoma|8251/3|BronchioloalveolarAdenocarcinoma
C739|ThyroidGland|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C739|ThyroidGland|826|PapillaryAdenocarcinoma|8260/3|PapillaryAdenocarcinoma
C739|ThyroidGland|826|PapillaryAdenocarcinoma|8261/2|AdenocarcinomaInSitu
C739|ThyroidGland|826|PapillaryAdenocarcinoma|8261/3|AdenocarcinomaInVillousAdenoma
C739|ThyroidGland|826|PapillaryAdenocarcinoma|8262/3|VillousAdenocarcinoma
C739|ThyroidGland|826|PapillaryAdenocarcinoma|8263/2|AdenocarcinomaInSitu
C739|ThyroidGland|826|PapillaryAdenocarcinoma|8263/3|AdenocarcinomaInTubulovillousAdenoma
C739|ThyroidGland|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C739|ThyroidGland|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C739|ThyroidGland|833|FollicularThyroidCarcinoma|8330/3|FollicularThyroidCarcinoma
C739|ThyroidGland|833|FollicularThyroidCarcinoma|8331/3|FollicularThyroidCarcinoma
C739|ThyroidGland|833|FollicularThyroidCarcinoma|8332/3|FollicularThyroidCarcinoma
C739|ThyroidGland|833|FollicularThyroidCarcinoma|8333/3|FetalAdenocarcinoma
C739|ThyroidGland|833|FollicularThyroidCarcinoma|8335/3|FollicularThyroidCarcinoma
C739|ThyroidGland|833|FollicularThyroidCarcinoma|8337/3|PoorlyDifferentiatedThyroidCarcinoma
C739|ThyroidGland|833|FollicularThyroidCarcinoma|8339/3|FollicularThyroidCarcinoma
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8340/3|PapillaryCarcinomaFollicularVariant
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8341/3|PapillaryMicrocarcinoma
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8342/3|PapillaryCarcinomaOxyphilicCell
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8343/2|PapillaryAndFollicularAdenocarcinoma
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8343/3|EncapsulatedPapillaryThyroidCarcinoma
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8344/3|PapillaryCarcinomaColumnarCell
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8345/3|MedullaryCarcinomaWithAmyloidStroma
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8346/3|MixedMedullaryfollicularCarcinoma
C739|ThyroidGland|834|PapillaryAndFollicularAdenocarcinoma|8347/3|MixedMedullarypapillaryCarcinoma
C739|ThyroidGland|835|NonencapsulatedSclerosingCarcinoma|8350/3|NonencapsulatedSclerosingCarcinoma
C739|ThyroidGland|845|PapillaryCystadenocarcinoma|8450/3|PapillaryCystadenocarcinoma
C739|ThyroidGland|851|MedullaryCarcinoma|8510/3|MedullaryCarcinoma
C739|ThyroidGland|855|AcinarCellCarcinoma|8550/3|AcinarCellCarcinoma
C739|ThyroidGland|855|AcinarCellCarcinoma|8551/3|AcinarCellCystadenocarcinoma
C739|ThyroidGland|883|BenignFibrousHistiocytoma|8830/3|MalignantFibrousHistiocytoma
C739|ThyroidGland|898|Carcinosarcoma|8980/3|Carcinosarcoma
C739|ThyroidGland|898|Carcinosarcoma|8981/3|CarcinosarcomaEmbryonal
C739|ThyroidGland|898|Carcinosarcoma|8982/3|MalignantMyoepithelioma
C739|ThyroidGland|959|Lymphoma|9590/3|Lymphoma
C739|ThyroidGland|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C739|ThyroidGland|959|Lymphoma|9596/3|CompositeLymphoma
C739|ThyroidGland|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C739|ThyroidGland|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C739|ThyroidGland|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C739|ThyroidGland|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C739|ThyroidGland|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C739|ThyroidGland|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C739|ThyroidGland|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C739|ThyroidGland|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C739|ThyroidGland|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C739|ThyroidGland|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C739|ThyroidGland|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C739|ThyroidGland|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C739|ThyroidGland|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C739|ThyroidGland|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C739|ThyroidGland|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C739|ThyroidGland|967|BCellLymphomas|9673/3|MantleCellLymphoma
C739|ThyroidGland|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C739|ThyroidGland|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C739|ThyroidGland|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C739|ThyroidGland|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C739|ThyroidGland|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C739|ThyroidGland|969|FollicularAdenoma|9690/3|LymphomaFollicular
C739|ThyroidGland|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C739|ThyroidGland|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C739|ThyroidGland|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C739|ThyroidGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C739|ThyroidGland|970|TCellLymphoma|9701/3|SezarySyndrome
C739|ThyroidGland|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C739|ThyroidGland|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C739|ThyroidGland|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C739|ThyroidGland|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C739|ThyroidGland|971|AdultNonHodgkinLymphoma|9715/3|AnaplasticLargeCellLymphoma
C739|ThyroidGland|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C739|ThyroidGland|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C739|ThyroidGland|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C739|ThyroidGland|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C739|ThyroidGland|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C739|ThyroidGland|973|Plasmacytoma|9731/3|Plasmacytoma
C739|ThyroidGland|973|Plasmacytoma|9734/3|ExtramedullaryPlasmacytoma
C739|ThyroidGland|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C739|ThyroidGland|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C739|ThyroidGland|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C739|ThyroidGland|974|MastCellNeoplasm|9740/3|MastCellSarcoma
C739|ThyroidGland|974|MastCellNeoplasm|9741/3|MalignantMastocytosis
C739|ThyroidGland|974|MastCellNeoplasm|9749/3|ErdheimChesterDisease
C739|ThyroidGland|975|TrueHistiocyticLymphoma|9750/3|MalignantHistiocytosis
C739|ThyroidGland|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C739|ThyroidGland|975|TrueHistiocyticLymphoma|9754/3|AdultLangerhansCellHistiocytosis
C739|ThyroidGland|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C739|ThyroidGland|975|TrueHistiocyticLymphoma|9756/3|LangerhansCellSarcoma
C739|ThyroidGland|975|TrueHistiocyticLymphoma|9757/3|InterdigitatingDendriticCellSarcoma
C739|ThyroidGland|975|TrueHistiocyticLymphoma|9758/3|FollicularDendriticCellSarcoma
C739|ThyroidGland|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C739|ThyroidGland|976|ImmunoproliferativeDisorder|9766/3|LymphomatoidGranulomatosis
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9812/3|null
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9813/3|null
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9814/3|null
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9817/3|null
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9818/3|null
C739|ThyroidGland|981|PrecursorLymphoidNeoplasm|9819/3|LeukemiaBCell
C739|ThyroidGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C739|ThyroidGland|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C739|ThyroidGland|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C739|ThyroidGland|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C739|ThyroidGland|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C739|ThyroidGland|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C739|ThyroidGland|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
C740-C741,C749|AdrenalGland|801|Carcinoma|8010/2|InSituCancer
C740-C741,C749|AdrenalGland|801|Carcinoma|8010/3|CarcinomaNOSDNE
C740-C741,C749|AdrenalGland|801|Carcinoma|8011/3|MalignantEpithelioma
C740-C741,C749|AdrenalGland|801|Carcinoma|8012/3|LargeCellCarcinoma
C740-C741,C749|AdrenalGland|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C740-C741,C749|AdrenalGland|801|Carcinoma|8014/3|LargeCellCarcinoma
C740-C741,C749|AdrenalGland|801|Carcinoma|8015/3|GlassyCellCarcinoma
C740-C741,C749|AdrenalGland|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C740-C741,C749|AdrenalGland|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C740-C741,C749|AdrenalGland|802|Carcinoma|8022/3|PleomorphicCarcinoma
C740-C741,C749|AdrenalGland|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C740-C741,C749|AdrenalGland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C740-C741,C749|AdrenalGland|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C740-C741,C749|AdrenalGland|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C740-C741,C749|AdrenalGland|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C740-C741,C749|AdrenalGland|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C740-C741,C749|AdrenalGland|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C740-C741,C749|AdrenalGland|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C740-C741,C749|AdrenalGland|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C740-C741,C749|AdrenalGland|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C740-C741,C749|AdrenalGland|837|AdrenocorticalCarcinoma|8370/3|AdrenocorticalCarcinoma
C740-C741,C749|AdrenalGland|868|Paraganglioma|8680/3|MalignantParaganglioma
C740-C741,C749|AdrenalGland|869|MalignantExtraAdrenalParaganglioma|8693/3|MalignantExtraAdrenalParaganglioma
C740-C741,C749|AdrenalGland|870|Pheochromocytoma|8700/3|Pheochromocytoma
C740-C741,C749|AdrenalGland|906|GermCellTumor|9060/3|Dysgerminoma
C740-C741,C749|AdrenalGland|906|GermCellTumor|9064/3|Germinoma
C740-C741,C749|AdrenalGland|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C740-C741,C749|AdrenalGland|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C740-C741,C749|AdrenalGland|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C740-C741,C749|AdrenalGland|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C740-C741,C749|AdrenalGland|908|Teratoma|9080/3|ImmatureTeratoma
C740-C741,C749|AdrenalGland|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C740-C741,C749|AdrenalGland|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C740-C741,C749|AdrenalGland|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C740-C741,C749|AdrenalGland|908|Teratoma|9084/3|Teratoma
C740-C741,C749|AdrenalGland|908|Teratoma|9085/3|MixedGermCellTumor
C740-C741,C749|AdrenalGland|937|Chordoma|9370/3|Chordoma
C740-C741,C749|AdrenalGland|937|Chordoma|9371/3|ChondroidChordoma
C740-C741,C749|AdrenalGland|937|Chordoma|9372/3|DedifferentiatedChordoma
C740-C741,C749|AdrenalGland|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C740-C741,C749|AdrenalGland|950|Neuroblastoma|9500/3|Neuroblastoma
C740-C741,C749|AdrenalGland|950|Neuroblastoma|9501/3|Medulloepithelioma
C740-C741,C749|AdrenalGland|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C740-C741,C749|AdrenalGland|950|Neuroblastoma|9503/3|Neuroepithelioma
C740-C741,C749|AdrenalGland|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C740-C741,C749|AdrenalGland|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C740-C741,C749|AdrenalGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C740-C741,C749|AdrenalGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C750|ParathyroidGland|801|Carcinoma|8010/2|InSituCancer
C750|ParathyroidGland|801|Carcinoma|8010/3|CarcinomaNOSDNE
C750|ParathyroidGland|801|Carcinoma|8011/3|MalignantEpithelioma
C750|ParathyroidGland|801|Carcinoma|8012/3|LargeCellCarcinoma
C750|ParathyroidGland|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C750|ParathyroidGland|801|Carcinoma|8014/3|LargeCellCarcinoma
C750|ParathyroidGland|801|Carcinoma|8015/3|GlassyCellCarcinoma
C750|ParathyroidGland|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C750|ParathyroidGland|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C750|ParathyroidGland|802|Carcinoma|8022/3|PleomorphicCarcinoma
C750|ParathyroidGland|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C750|ParathyroidGland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C750|ParathyroidGland|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C750|ParathyroidGland|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C750|ParathyroidGland|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C750|ParathyroidGland|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C750|ParathyroidGland|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C750|ParathyroidGland|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C750|ParathyroidGland|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C750|ParathyroidGland|832|GranularCellCarcinoma|8322/3|WaterClearCellAdenocarcinoma
C750|ParathyroidGland|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C750|ParathyroidGland|868|Paraganglioma|8680/3|MalignantParaganglioma
C750|ParathyroidGland|869|MalignantExtraAdrenalParaganglioma|8693/3|MalignantExtraAdrenalParaganglioma
C750|ParathyroidGland|906|GermCellTumor|9060/3|Dysgerminoma
C750|ParathyroidGland|906|GermCellTumor|9064/3|Germinoma
C750|ParathyroidGland|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C750|ParathyroidGland|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C750|ParathyroidGland|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C750|ParathyroidGland|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C750|ParathyroidGland|908|Teratoma|9080/3|ImmatureTeratoma
C750|ParathyroidGland|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C750|ParathyroidGland|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C750|ParathyroidGland|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C750|ParathyroidGland|908|Teratoma|9084/3|Teratoma
C750|ParathyroidGland|908|Teratoma|9085/3|MixedGermCellTumor
C750|ParathyroidGland|937|Chordoma|9370/3|Chordoma
C750|ParathyroidGland|937|Chordoma|9371/3|ChondroidChordoma
C750|ParathyroidGland|937|Chordoma|9372/3|DedifferentiatedChordoma
C750|ParathyroidGland|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C750|ParathyroidGland|950|Neuroblastoma|9500/3|Neuroblastoma
C750|ParathyroidGland|950|Neuroblastoma|9501/3|Medulloepithelioma
C750|ParathyroidGland|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C750|ParathyroidGland|950|Neuroblastoma|9503/3|Neuroepithelioma
C750|ParathyroidGland|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C750|ParathyroidGland|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C750|ParathyroidGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C750|ParathyroidGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C751|PituitaryGland|801|Carcinoma|8010/0|BenignEpithelioma
C751|PituitaryGland|801|Carcinoma|8010/2|InSituCancer
C751|PituitaryGland|801|Carcinoma|8010/3|CarcinomaNOSDNE
C751|PituitaryGland|814|Adenocarcinoma|8140/0|Adenoma
C751|PituitaryGland|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C751|PituitaryGland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C751|PituitaryGland|814|Adenocarcinoma|8146/0|SalivaryGlandMonomorphicAdenoma
C751|PituitaryGland|826|PapillaryAdenocarcinoma|8260/0|PapillaryAdenoma
C751|PituitaryGland|827|ChromophobeRenalCellCarcinoma|8270/0|PituitaryGlandChromophobeAdenoma
C751|PituitaryGland|827|ChromophobeRenalCellCarcinoma|8270/3|ChromophobeRenalCellCarcinoma
C751|PituitaryGland|827|ChromophobeRenalCellCarcinoma|8271/0|Prolactinoma
C751|PituitaryGland|827|ChromophobeRenalCellCarcinoma|8272/0|PituitaryAdenoma
C751|PituitaryGland|827|ChromophobeRenalCellCarcinoma|8272/3|PituitaryCarcinoma
C751|PituitaryGland|827|ChromophobeRenalCellCarcinoma|8273/3|Blastoma
C751|PituitaryGland|828|AcidophilCarcinoma|8280/0|PituitaryGlandAcidophilAdenoma
C751|PituitaryGland|828|AcidophilCarcinoma|8280/3|AcidophilCarcinoma
C751|PituitaryGland|828|AcidophilCarcinoma|8281/0|MixedAcidophilbasophilAdenoma
C751|PituitaryGland|828|AcidophilCarcinoma|8281/3|MixedAcidophilbasophilCarcinoma
C751|PituitaryGland|829|OxyphilicAdenocarcinoma|8290/0|OxyphilicAdenoma
C751|PituitaryGland|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C751|PituitaryGland|830|BasophilicAdenocarcinoma|8300/0|PituitaryGlandBasophilAdenoma
C751|PituitaryGland|830|BasophilicAdenocarcinoma|8300/3|BasophilicAdenocarcinoma
C751|PituitaryGland|831|ClearCellAdenocarcinoma|8310/0|ClearCellAdenoma
C751|PituitaryGland|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C751|PituitaryGland|832|GranularCellCarcinoma|8323/0|MixedCellAdenoma
C751|PituitaryGland|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C751|PituitaryGland|880|Sarcoma|8800/0|BenignSoftTissueNeoplasm
C751|PituitaryGland|880|Sarcoma|8800/3|Sarcoma
C751|PituitaryGland|885|Liposarcoma|8850/0|Lipoma
C751|PituitaryGland|906|GermCellTumor|9060/3|Dysgerminoma
C751|PituitaryGland|906|GermCellTumor|9064/3|Germinoma
C751|PituitaryGland|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C751|PituitaryGland|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C751|PituitaryGland|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C751|PituitaryGland|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C751|PituitaryGland|908|Teratoma|9080/0|MatureTeratoma
C751|PituitaryGland|908|Teratoma|9080/1|Teratoma
C751|PituitaryGland|908|Teratoma|9080/3|ImmatureTeratoma
C751|PituitaryGland|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C751|PituitaryGland|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C751|PituitaryGland|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C751|PituitaryGland|908|Teratoma|9084/3|Teratoma
C751|PituitaryGland|908|Teratoma|9085/3|MixedGermCellTumor
C751|PituitaryGland|935|Craniopharyngioma|9350/1|Craniopharyngioma
C751|PituitaryGland|935|Craniopharyngioma|9351/1|AdamantinousCraniopharyngioma
C751|PituitaryGland|935|Craniopharyngioma|9352/1|PapillaryCraniopharyngioma
C751|PituitaryGland|937|Chordoma|9370/3|Chordoma
C751|PituitaryGland|937|Chordoma|9371/3|ChondroidChordoma
C751|PituitaryGland|937|Chordoma|9372/3|DedifferentiatedChordoma
C751|PituitaryGland|943|Astroblastoma|9432/1|Pituicytoma
C751|PituitaryGland|950|Neuroblastoma|9500/3|Neuroblastoma
C751|PituitaryGland|950|Neuroblastoma|9501/3|Medulloepithelioma
C751|PituitaryGland|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C751|PituitaryGland|950|Neuroblastoma|9503/3|Neuroepithelioma
C751|PituitaryGland|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C751|PituitaryGland|958|GranularCellTumor|9580/0|GranularCellTumor
C751|PituitaryGland|958|GranularCellTumor|9582/0|GranularCellTumor
C751|PituitaryGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C751|PituitaryGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C752|CraniopharyngealDuct|801|Carcinoma|8010/0|BenignEpithelioma
C752|CraniopharyngealDuct|801|Carcinoma|8010/2|InSituCancer
C752|CraniopharyngealDuct|801|Carcinoma|8010/3|CarcinomaNOSDNE
C752|CraniopharyngealDuct|814|Adenocarcinoma|8140/0|Adenoma
C752|CraniopharyngealDuct|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C752|CraniopharyngealDuct|814|Adenocarcinoma|8140/3|Adenocarcinoma
C752|CraniopharyngealDuct|814|Adenocarcinoma|8146/0|SalivaryGlandMonomorphicAdenoma
C752|CraniopharyngealDuct|826|PapillaryAdenocarcinoma|8260/0|PapillaryAdenoma
C752|CraniopharyngealDuct|827|ChromophobeRenalCellCarcinoma|8270/0|PituitaryGlandChromophobeAdenoma
C752|CraniopharyngealDuct|827|ChromophobeRenalCellCarcinoma|8270/3|ChromophobeRenalCellCarcinoma
C752|CraniopharyngealDuct|827|ChromophobeRenalCellCarcinoma|8271/0|Prolactinoma
C752|CraniopharyngealDuct|827|ChromophobeRenalCellCarcinoma|8272/0|PituitaryAdenoma
C752|CraniopharyngealDuct|827|ChromophobeRenalCellCarcinoma|8272/3|PituitaryCarcinoma
C752|CraniopharyngealDuct|828|AcidophilCarcinoma|8280/0|PituitaryGlandAcidophilAdenoma
C752|CraniopharyngealDuct|828|AcidophilCarcinoma|8280/3|AcidophilCarcinoma
C752|CraniopharyngealDuct|828|AcidophilCarcinoma|8281/0|MixedAcidophilbasophilAdenoma
C752|CraniopharyngealDuct|828|AcidophilCarcinoma|8281/3|MixedAcidophilbasophilCarcinoma
C752|CraniopharyngealDuct|829|OxyphilicAdenocarcinoma|8290/0|OxyphilicAdenoma
C752|CraniopharyngealDuct|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C752|CraniopharyngealDuct|830|BasophilicAdenocarcinoma|8300/0|PituitaryGlandBasophilAdenoma
C752|CraniopharyngealDuct|830|BasophilicAdenocarcinoma|8300/3|BasophilicAdenocarcinoma
C752|CraniopharyngealDuct|831|ClearCellAdenocarcinoma|8310/0|ClearCellAdenoma
C752|CraniopharyngealDuct|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C752|CraniopharyngealDuct|832|GranularCellCarcinoma|8323/0|MixedCellAdenoma
C752|CraniopharyngealDuct|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C752|CraniopharyngealDuct|880|Sarcoma|8800/0|BenignSoftTissueNeoplasm
C752|CraniopharyngealDuct|880|Sarcoma|8800/3|Sarcoma
C752|CraniopharyngealDuct|885|Liposarcoma|8850/0|Lipoma
C752|CraniopharyngealDuct|906|GermCellTumor|9060/3|Dysgerminoma
C752|CraniopharyngealDuct|906|GermCellTumor|9064/3|Germinoma
C752|CraniopharyngealDuct|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C752|CraniopharyngealDuct|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C752|CraniopharyngealDuct|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C752|CraniopharyngealDuct|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C752|CraniopharyngealDuct|908|Teratoma|9080/0|MatureTeratoma
C752|CraniopharyngealDuct|908|Teratoma|9080/1|Teratoma
C752|CraniopharyngealDuct|908|Teratoma|9080/3|ImmatureTeratoma
C752|CraniopharyngealDuct|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C752|CraniopharyngealDuct|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C752|CraniopharyngealDuct|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C752|CraniopharyngealDuct|908|Teratoma|9084/3|Teratoma
C752|CraniopharyngealDuct|908|Teratoma|9085/3|MixedGermCellTumor
C752|CraniopharyngealDuct|935|Craniopharyngioma|9350/1|Craniopharyngioma
C752|CraniopharyngealDuct|935|Craniopharyngioma|9351/1|AdamantinousCraniopharyngioma
C752|CraniopharyngealDuct|935|Craniopharyngioma|9352/1|PapillaryCraniopharyngioma
C752|CraniopharyngealDuct|937|Chordoma|9370/3|Chordoma
C752|CraniopharyngealDuct|937|Chordoma|9371/3|ChondroidChordoma
C752|CraniopharyngealDuct|937|Chordoma|9372/3|DedifferentiatedChordoma
C752|CraniopharyngealDuct|950|Neuroblastoma|9500/3|Neuroblastoma
C752|CraniopharyngealDuct|950|Neuroblastoma|9501/3|Medulloepithelioma
C752|CraniopharyngealDuct|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C752|CraniopharyngealDuct|950|Neuroblastoma|9503/3|Neuroepithelioma
C752|CraniopharyngealDuct|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C752|CraniopharyngealDuct|958|GranularCellTumor|9580/0|GranularCellTumor
C752|CraniopharyngealDuct|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C752|CraniopharyngealDuct|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C753|PinealGland|801|Carcinoma|8010/0|BenignEpithelioma
C753|PinealGland|906|GermCellTumor|9060/3|Dysgerminoma
C753|PinealGland|906|GermCellTumor|9064/3|Germinoma
C753|PinealGland|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C753|PinealGland|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C753|PinealGland|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C753|PinealGland|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C753|PinealGland|908|Teratoma|9080/0|MatureTeratoma
C753|PinealGland|908|Teratoma|9080/3|ImmatureTeratoma
C753|PinealGland|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C753|PinealGland|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C753|PinealGland|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C753|PinealGland|908|Teratoma|9084/0|DermoidCyst
C753|PinealGland|908|Teratoma|9084/3|Teratoma
C753|PinealGland|908|Teratoma|9085/3|MixedGermCellTumor
C753|PinealGland|936|NeuroepitheliomaPeripheral|9360/1|PinealGlandNeoplasm
C753|PinealGland|936|NeuroepitheliomaPeripheral|9361/1|Pineocytoma
C753|PinealGland|936|NeuroepitheliomaPeripheral|9362/3|Pineoblastoma
C753|PinealGland|937|Chordoma|9370/3|Chordoma
C753|PinealGland|937|Chordoma|9371/3|ChondroidChordoma
C753|PinealGland|937|Chordoma|9372/3|DedifferentiatedChordoma
C753|PinealGland|939|Ependymoma|9395/3|TumorOfThePinealRegion
C753|PinealGland|947|Medulloblastoma|9473/3|PrimitiveNeuroectodermalTumor
C753|PinealGland|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C753|PinealGland|949|Ganglioneuroblastoma|9492/0|Gangliocytoma
C753|PinealGland|950|Neuroblastoma|9500/3|Neuroblastoma
C753|PinealGland|950|Neuroblastoma|9501/3|Medulloepithelioma
C753|PinealGland|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C753|PinealGland|950|Neuroblastoma|9503/3|Neuroepithelioma
C753|PinealGland|950|Neuroblastoma|9505/1|Ganglioglioma
C753|PinealGland|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C753|PinealGland|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C753|PinealGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C753|PinealGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C754-C755,C758-C759|EndocrineGland|801|Carcinoma|8010/2|InSituCancer
C754-C755,C758-C759|EndocrineGland|801|Carcinoma|8010/3|CarcinomaNOSDNE
C754-C755,C758-C759|EndocrineGland|801|Carcinoma|8011/3|MalignantEpithelioma
C754-C755,C758-C759|EndocrineGland|801|Carcinoma|8012/3|LargeCellCarcinoma
C754-C755,C758-C759|EndocrineGland|801|Carcinoma|8013/3|LargeCellNeuroendocrineCarcinoma
C754-C755,C758-C759|EndocrineGland|801|Carcinoma|8014/3|LargeCellCarcinoma
C754-C755,C758-C759|EndocrineGland|801|Carcinoma|8015/3|GlassyCellCarcinoma
C754-C755,C758-C759|EndocrineGland|802|Carcinoma|8020/3|UndifferentiatedCarcinoma
C754-C755,C758-C759|EndocrineGland|802|Carcinoma|8021/3|AnaplasticCarcinomaDNE
C754-C755,C758-C759|EndocrineGland|802|Carcinoma|8022/3|PleomorphicCarcinoma
C754-C755,C758-C759|EndocrineGland|814|Adenocarcinoma|8140/2|AdenocarcinomaInSitu
C754-C755,C758-C759|EndocrineGland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C754-C755,C758-C759|EndocrineGland|814|Adenocarcinoma|8141/3|ScirrhousAdenocarcinoma
C754-C755,C758-C759|EndocrineGland|814|Adenocarcinoma|8143/3|SuperficialSpreadingAdenocarcinoma
C754-C755,C758-C759|EndocrineGland|814|Adenocarcinoma|8147/3|AdenocarcinomaBasalCell
C754-C755,C758-C759|EndocrineGland|825|BronchioloalveolarAdenocarcinoma|8255/3|AdenocarcinomaWithMixedSubtypes
C754-C755,C758-C759|EndocrineGland|829|OxyphilicAdenocarcinoma|8290/3|OxyphilicAdenocarcinoma
C754-C755,C758-C759|EndocrineGland|831|ClearCellAdenocarcinoma|8310/3|ClearCellAdenocarcinoma
C754-C755,C758-C759|EndocrineGland|832|GranularCellCarcinoma|8320/3|GranularCellCarcinoma
C754-C755,C758-C759|EndocrineGland|832|GranularCellCarcinoma|8323/3|MixedCellAdenocarcinoma
C754-C755,C758-C759|EndocrineGland|868|Paraganglioma|8680/3|MalignantParaganglioma
C754-C755,C758-C759|EndocrineGland|868|Paraganglioma|8681/3|SympatheticParaganglioma
C754-C755,C758-C759|EndocrineGland|868|Paraganglioma|8682/3|ParasympatheticParaganglioma
C754-C755,C758-C759|EndocrineGland|869|MalignantExtraAdrenalParaganglioma|8690/3|MiddleEarParaganglioma
C754-C755,C758-C759|EndocrineGland|869|MalignantExtraAdrenalParaganglioma|8691/3|AorticopulmonaryParaganglioma
C754-C755,C758-C759|EndocrineGland|869|MalignantExtraAdrenalParaganglioma|8692/3|CarotidBodyParaganglioma
C754-C755,C758-C759|EndocrineGland|869|MalignantExtraAdrenalParaganglioma|8693/3|MalignantExtraAdrenalParaganglioma
C754-C755,C758-C759|EndocrineGland|906|GermCellTumor|9060/3|Dysgerminoma
C754-C755,C758-C759|EndocrineGland|906|GermCellTumor|9064/3|Germinoma
C754-C755,C758-C759|EndocrineGland|906|GermCellTumor|9065/3|NongerminomatousGermCellTumorC1266158
C754-C755,C758-C759|EndocrineGland|907|EmbryonalCarcinoma|9070/3|EmbryonalCarcinoma
C754-C755,C758-C759|EndocrineGland|907|EmbryonalCarcinoma|9071/3|YolkSacTumor
C754-C755,C758-C759|EndocrineGland|907|EmbryonalCarcinoma|9072/3|Polyembryoma
C754-C755,C758-C759|EndocrineGland|908|Teratoma|9080/3|ImmatureTeratoma
C754-C755,C758-C759|EndocrineGland|908|Teratoma|9081/3|MixedEmbryonalCarcinomaAndTeratoma
C754-C755,C758-C759|EndocrineGland|908|Teratoma|9082/3|UndifferentiatedImmatureTeratoma
C754-C755,C758-C759|EndocrineGland|908|Teratoma|9083/3|IntermediateImmatureTeratoma
C754-C755,C758-C759|EndocrineGland|908|Teratoma|9084/3|Teratoma
C754-C755,C758-C759|EndocrineGland|908|Teratoma|9085/3|MixedGermCellTumor
C754-C755,C758-C759|EndocrineGland|937|Chordoma|9370/3|Chordoma
C754-C755,C758-C759|EndocrineGland|937|Chordoma|9371/3|ChondroidChordoma
C754-C755,C758-C759|EndocrineGland|937|Chordoma|9372/3|DedifferentiatedChordoma
C754-C755,C758-C759|EndocrineGland|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C754-C755,C758-C759|EndocrineGland|950|Neuroblastoma|9500/3|Neuroblastoma
C754-C755,C758-C759|EndocrineGland|950|Neuroblastoma|9501/3|Medulloepithelioma
C754-C755,C758-C759|EndocrineGland|950|Neuroblastoma|9502/3|TeratoidMedulloepithelioma
C754-C755,C758-C759|EndocrineGland|950|Neuroblastoma|9503/3|Neuroepithelioma
C754-C755,C758-C759|EndocrineGland|950|Neuroblastoma|9504/3|PolarSpongioblastoma
C754-C755,C758-C759|EndocrineGland|950|Neuroblastoma|9505/3|AnaplasticGanglioglioma
C754-C755,C758-C759|EndocrineGland|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C754-C755,C758-C759|EndocrineGland|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C770-C775,C778-C779|LymphNode|959|Lymphoma|9590/3|Lymphoma
C770-C775,C778-C779|LymphNode|959|Lymphoma|9591/3|AdultNonHodgkinLymphoma
C770-C775,C778-C779|LymphNode|959|Lymphoma|9596/3|CompositeLymphoma
C770-C775,C778-C779|LymphNode|965|AdultHodgkinLymphoma|9650/3|AdultHodgkinLymphoma
C770-C775,C778-C779|LymphNode|965|AdultHodgkinLymphoma|9651/3|HodgkinLymphomaLymphocyterich
C770-C775,C778-C779|LymphNode|965|AdultHodgkinLymphoma|9652/3|MixedCellularityHodgkinLymphoma
C770-C775,C778-C779|LymphNode|965|AdultHodgkinLymphoma|9653/3|ChronicLymphocyticLeukemia
C770-C775,C778-C779|LymphNode|965|AdultHodgkinLymphoma|9654/3|HodgkinLymphomaLymphocyteDepletion
C770-C775,C778-C779|LymphNode|965|AdultHodgkinLymphoma|9655/3|AdultHodgkinLymphoma
C770-C775,C778-C779|LymphNode|965|AdultHodgkinLymphoma|9659/3|ChildhoodNLPHD
C770-C775,C778-C779|LymphNode|966|AdultHodgkinLymphoma|9661/3|HodgkinsGranuloma
C770-C775,C778-C779|LymphNode|966|AdultHodgkinLymphoma|9662/3|HodgkinSarcomaObsolete
C770-C775,C778-C779|LymphNode|966|AdultHodgkinLymphoma|9663/3|HodgkinsNodularSclerosis
C770-C775,C778-C779|LymphNode|966|AdultHodgkinLymphoma|9664/3|HodgkinSclerCellDNE
C770-C775,C778-C779|LymphNode|966|AdultHodgkinLymphoma|9665/3|HodgkinLymphomaGrade1DNE
C770-C775,C778-C779|LymphNode|966|AdultHodgkinLymphoma|9667/3|HodgkinLymphomaGrade2DNE
C770-C775,C778-C779|LymphNode|967|BCellLymphomas|9670/3|SmallLymphocyticLymphoma
C770-C775,C778-C779|LymphNode|967|BCellLymphomas|9671/3|LymphoplasmacyticLymphoma
C770-C775,C778-C779|LymphNode|967|BCellLymphomas|9673/3|MantleCellLymphoma
C770-C775,C778-C779|LymphNode|967|BCellLymphomas|9675/3|DiffuseMalignantLymphoma
C770-C775,C778-C779|LymphNode|967|BCellLymphomas|9678/3|PrimaryEffusionLymphoma
C770-C775,C778-C779|LymphNode|967|BCellLymphomas|9679/3|MediastinalLargeBcellLymphoma
C770-C775,C778-C779|LymphNode|968|DiffuseLargeBCellLymphoma|9680/3|DiffuseLargeBCellLymphoma
C770-C775,C778-C779|LymphNode|968|DiffuseLargeBCellLymphoma|9684/3|ImmunoblasticLymphoma
C770-C775,C778-C779|LymphNode|968|DiffuseLargeBCellLymphoma|9687/3|BurkittLymphoma
C770-C775,C778-C779|LymphNode|968|DiffuseLargeBCellLymphoma|9688/3|BCellNonHodgkinLymphoma
C770-C775,C778-C779|LymphNode|968|DiffuseLargeBCellLymphoma|9689/3|MucosaassociatedLymphoma
C770-C775,C778-C779|LymphNode|969|FollicularAdenoma|9690/3|LymphomaFollicular
C770-C775,C778-C779|LymphNode|969|FollicularAdenoma|9691/3|Grade2FollicularLymphoma
C770-C775,C778-C779|LymphNode|969|FollicularAdenoma|9695/3|FollicularLymphomaGrade1
C770-C775,C778-C779|LymphNode|969|FollicularAdenoma|9698/3|LymphomaFollicularGrade3
C770-C775,C778-C779|LymphNode|969|FollicularAdenoma|9699/3|MucosaassociatedLymphoma
C770-C775,C778-C779|LymphNode|970|TCellLymphoma|9702/3|PeripheralTCellLymphoma
C770-C775,C778-C779|LymphNode|970|TCellLymphoma|9705/3|AngioimmunoblasticLymphadenopathy
C770-C775,C778-C779|LymphNode|970|TCellLymphoma|9708/3|TCellLymphoma
C770-C775,C778-C779|LymphNode|971|AdultNonHodgkinLymphoma|9712/3|Angioendotheliomatosis
C770-C775,C778-C779|LymphNode|971|AdultNonHodgkinLymphoma|9714/3|AnaplasticLargeCellLymphoma
C770-C775,C778-C779|LymphNode|971|AdultNonHodgkinLymphoma|9716/3|Lymphoma
C770-C775,C778-C779|LymphNode|971|AdultNonHodgkinLymphoma|9717/3|IntestinalTCellLymphomaNOS
C770-C775,C778-C779|LymphNode|971|AdultNonHodgkinLymphoma|9719/3|TCellLymphoma
C770-C775,C778-C779|LymphNode|972|LymphoblasticLymphoma|9724/3|LymphoproliferativeDisorder
C770-C775,C778-C779|LymphNode|972|LymphoblasticLymphoma|9727/3|LymphoblasticLymphoma
C770-C775,C778-C779|LymphNode|972|LymphoblasticLymphoma|9728/3|PrecursorBLymphoblast
C770-C775,C778-C779|LymphNode|972|LymphoblasticLymphoma|9729/3|PrecursorTLymphoblast
C770-C775,C778-C779|LymphNode|973|Plasmacytoma|9735/3|PlasmablasticLymphoma
C770-C775,C778-C779|LymphNode|973|Plasmacytoma|9737/3|BCellNonHodgkinLymphoma
C770-C775,C778-C779|LymphNode|973|Plasmacytoma|9738/3|BCellNonHodgkinLymphomaDNE
C770-C775,C778-C779|LymphNode|975|TrueHistiocyticLymphoma|9751/3|AdultLangerhansCellHistiocytosis
C770-C775,C778-C779|LymphNode|975|TrueHistiocyticLymphoma|9755/3|HistiocyticSarcoma
C770-C775,C778-C779|LymphNode|975|TrueHistiocyticLymphoma|9759/3|FibroblasticReticularCellTumor
C770-C775,C778-C779|LymphNode|976|ImmunoproliferativeDisorder|9761/3|WaldenstromMacroglobulinemia
C770-C775,C778-C779|LymphNode|976|ImmunoproliferativeDisorder|9762/3|HeavyChainDisease
C770-C775,C778-C779|LymphNode|981|PrecursorLymphoidNeoplasm|9811/3|BLymphoblasticLeukemiaLymphoma
C770-C775,C778-C779|LymphNode|981|PrecursorLymphoidNeoplasm|9812/3|null
C770-C775,C778-C779|LymphNode|981|PrecursorLymphoidNeoplasm|9813/3|null
C770-C775,C778-C779|LymphNode|981|PrecursorLymphoidNeoplasm|9814/3|null
C770-C775,C778-C779|LymphNode|981|PrecursorLymphoidNeoplasm|9815/3|BLymphoblasticLeukemiaLymphoma
C770-C775,C778-C779|LymphNode|981|PrecursorLymphoidNeoplasm|9816/3|HypodiploidALL
C770-C775,C778-C779|LymphNode|981|PrecursorLymphoidNeoplasm|9817/3|null
C770-C775,C778-C779|LymphNode|981|PrecursorLymphoidNeoplasm|9818/3|null
C770-C775,C778-C779|LymphNode|982|LymphoidLeukemia|9823/3|ChronicLymphocyticLeukemia
C770-C775,C778-C779|LymphNode|983|Leukemia|9831/3|LeukemiaLargeGranularLymphocytic
C770-C775,C778-C779|LymphNode|983|Leukemia|9837/3|TLymphoblasticLeukemiaLymphoma
C770-C775,C778-C779|LymphNode|996|MyeloproliferativeNeoplasm|9965/3|LymphocyticNeoplasm
C770-C775,C778-C779|LymphNode|996|MyeloproliferativeNeoplasm|9967/3|LymphocyticNeoplasm
C770-C775,C778-C779|LymphNode|997|MyeloproliferativeNeoplasm|9971/3|PolymorphicPTLD
C770-C775,C778-C779|LymphNode|997|MyeloproliferativeNeoplasm|9975/3|MyeloproliferativeNeoplasm
