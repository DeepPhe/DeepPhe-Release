-cancer ID|*patient ID|*body location|body location laterality|Temporality|clinical stage|clinical T classification|clinical N classification|clinical M classification|-clinical prefix|-clinical suffix|pathologic T classification|pathologic N classification|pathologic M classification|-pathologic prefix|-pathologic suffixcancer_patientX_Left_Breast_Current|patientX|Breast|Left|Current|Stage_2A|cT1_Stage_Finding|cN1_Stage_Finding|cM0_Stage_Finding|||pT1c_Stage_Finding|pN1a_Stage_Finding|||