C000-C006,C008-C009|Lip_Proper|800|Neoplasm|8000/3|Malignant_Neoplasm
C000-C006,C008-C009|Lip_Proper|800|Neoplasm|8001/3|Malignant_Cell
C000-C006,C008-C009|Lip_Proper|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C000-C006,C008-C009|Lip_Proper|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C000-C006,C008-C009|Lip_Proper|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C000-C006,C008-C009|Lip_Proper|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C000-C006,C008-C009|Lip_Proper|801|Carcinoma|8010/2|In_Situ_Cancer
C000-C006,C008-C009|Lip_Proper|801|Carcinoma|8010/3|Carcinoma
C000-C006,C008-C009|Lip_Proper|801|Carcinoma|8011/3|Malignant_Epithelioma
C000-C006,C008-C009|Lip_Proper|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C000-C006,C008-C009|Lip_Proper|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C000-C006,C008-C009|Lip_Proper|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C000-C006,C008-C009|Lip_Proper|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C000-C006,C008-C009|Lip_Proper|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C000-C006,C008-C009|Lip_Proper|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C000-C006,C008-C009|Lip_Proper|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C000-C006,C008-C009|Lip_Proper|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C000-C006,C008-C009|Lip_Proper|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C000-C006,C008-C009|Lip_Proper|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C000-C006,C008-C009|Lip_Proper|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C000-C006,C008-C009|Lip_Proper|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C000-C006,C008-C009|Lip_Proper|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C000-C006,C008-C009|Lip_Proper|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C000-C006,C008-C009|Lip_Proper|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C000-C006,C008-C009|Lip_Proper|814|Adenocarcinoma|8140/3|Adenocarcinoma
C000-C006,C008-C009|Lip_Proper|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C000-C006,C008-C009|Lip_Proper|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C000-C006,C008-C009|Lip_Proper|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C000-C006,C008-C009|Lip_Proper|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C000-C006,C008-C009|Lip_Proper|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C000-C006,C008-C009|Lip_Proper|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C000-C006,C008-C009|Lip_Proper|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C000-C006,C008-C009|Lip_Proper|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C000-C006,C008-C009|Lip_Proper|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C000-C006,C008-C009|Lip_Proper|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C000-C006,C008-C009|Lip_Proper|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C000-C006,C008-C009|Lip_Proper|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C000-C006,C008-C009|Lip_Proper|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C000-C006,C008-C009|Lip_Proper|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C000-C006,C008-C009|Lip_Proper|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C000-C006,C008-C009|Lip_Proper|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C000-C006,C008-C009|Lip_Proper|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C000-C006,C008-C009|Lip_Proper|872|Melanoma|8720/3|Melanoma
C000-C006,C008-C009|Lip_Proper|872|Melanoma|8721/3|Nodular_Melanoma
C000-C006,C008-C009|Lip_Proper|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C000-C006,C008-C009|Lip_Proper|872|Melanoma|8723/3|Regressing_Melanoma
C000-C006,C008-C009|Lip_Proper|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C000-C006,C008-C009|Lip_Proper|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C000-C006,C008-C009|Lip_Proper|874|Nevus|8745/3|Desmoplastic_Melanoma
C000-C006,C008-C009|Lip_Proper|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C000-C006,C008-C009|Lip_Proper|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C000-C006,C008-C009|Lip_Proper|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C000-C006,C008-C009|Lip_Proper|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C000-C006,C008-C009|Lip_Proper|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C000-C006,C008-C009|Lip_Proper|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C000-C006,C008-C009|Lip_Proper|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C000-C006,C008-C009|Lip_Proper|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C000-C006,C008-C009|Lip_Proper|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C019|Root_Of_Tongue|800|Neoplasm|8000/3|Malignant_Neoplasm
C019|Root_Of_Tongue|800|Neoplasm|8001/3|Malignant_Cell
C019|Root_Of_Tongue|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C019|Root_Of_Tongue|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C019|Root_Of_Tongue|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C019|Root_Of_Tongue|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C019|Root_Of_Tongue|801|Carcinoma|8010/2|In_Situ_Cancer
C019|Root_Of_Tongue|801|Carcinoma|8010/3|Carcinoma
C019|Root_Of_Tongue|801|Carcinoma|8011/3|Malignant_Epithelioma
C019|Root_Of_Tongue|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C019|Root_Of_Tongue|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C019|Root_Of_Tongue|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C019|Root_Of_Tongue|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C019|Root_Of_Tongue|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C019|Root_Of_Tongue|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C019|Root_Of_Tongue|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C019|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C019|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C019|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C019|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C019|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C019|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C019|Root_Of_Tongue|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C019|Root_Of_Tongue|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C019|Root_Of_Tongue|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C019|Root_Of_Tongue|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C019|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C019|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C019|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8085/3|Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8086/3|Squamous_Cell_Carcinoma
C019|Root_Of_Tongue|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C019|Root_Of_Tongue|814|Adenocarcinoma|8140/3|Adenocarcinoma
C019|Root_Of_Tongue|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C019|Root_Of_Tongue|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C019|Root_Of_Tongue|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C019|Root_Of_Tongue|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C019|Root_Of_Tongue|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C019|Root_Of_Tongue|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C019|Root_Of_Tongue|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C019|Root_Of_Tongue|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C019|Root_Of_Tongue|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C019|Root_Of_Tongue|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C019|Root_Of_Tongue|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C019|Root_Of_Tongue|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C019|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C019|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C019|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C019|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C019|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C019|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C019|Root_Of_Tongue|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C019|Root_Of_Tongue|872|Melanoma|8720/3|Melanoma
C019|Root_Of_Tongue|872|Melanoma|8721/3|Nodular_Melanoma
C019|Root_Of_Tongue|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C019|Root_Of_Tongue|872|Melanoma|8723/3|Regressing_Melanoma
C019|Root_Of_Tongue|882|Sarcoma|8825/3|Sarcoma
C019|Root_Of_Tongue|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C019|Root_Of_Tongue|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C019|Root_Of_Tongue|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C019|Root_Of_Tongue|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C019|Root_Of_Tongue|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C019|Root_Of_Tongue|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C019|Root_Of_Tongue|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C019|Root_Of_Tongue|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C019|Root_Of_Tongue|959|Lymphoma|9590/3|Lymphoma
C019|Root_Of_Tongue|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C019|Root_Of_Tongue|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C019|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C019|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C019|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C019|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C019|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C019|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C019|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C019|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C019|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C019|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C019|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C019|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C019|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C019|Root_Of_Tongue|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C019|Root_Of_Tongue|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C019|Root_Of_Tongue|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C019|Root_Of_Tongue|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C019|Root_Of_Tongue|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C019|Root_Of_Tongue|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C019|Root_Of_Tongue|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C019|Root_Of_Tongue|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C019|Root_Of_Tongue|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C019|Root_Of_Tongue|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C019|Root_Of_Tongue|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C019|Root_Of_Tongue|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C019|Root_Of_Tongue|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C019|Root_Of_Tongue|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C019|Root_Of_Tongue|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C019|Root_Of_Tongue|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C019|Root_Of_Tongue|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C019|Root_Of_Tongue|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C019|Root_Of_Tongue|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C019|Root_Of_Tongue|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C019|Root_Of_Tongue|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C019|Root_Of_Tongue|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C019|Root_Of_Tongue|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C019|Root_Of_Tongue|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C019|Root_Of_Tongue|973|Plasmacytoma|9731/3|Plasmacytoma
C019|Root_Of_Tongue|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C019|Root_Of_Tongue|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C019|Root_Of_Tongue|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C019|Root_Of_Tongue|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C019|Root_Of_Tongue|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C019|Root_Of_Tongue|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C019|Root_Of_Tongue|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C019|Root_Of_Tongue|975|Neoplasm|9750/3|Malignant_Histiocytosis
C019|Root_Of_Tongue|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C019|Root_Of_Tongue|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C019|Root_Of_Tongue|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C019|Root_Of_Tongue|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C019|Root_Of_Tongue|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C019|Root_Of_Tongue|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C019|Root_Of_Tongue|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C019|Root_Of_Tongue|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C019|Root_Of_Tongue|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C019|Root_Of_Tongue|981|Neoplasm|9812/3|Lymphoma
C019|Root_Of_Tongue|981|Neoplasm|9813/3|Lymphoma
C019|Root_Of_Tongue|981|Neoplasm|9814/3|Lymphoma
C019|Root_Of_Tongue|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C019|Root_Of_Tongue|981|Neoplasm|9816/3|Hypodiploid_ALL
C019|Root_Of_Tongue|981|Neoplasm|9817/3|Lymphoma
C019|Root_Of_Tongue|981|Neoplasm|9818/3|Lymphoma
C019|Root_Of_Tongue|981|Neoplasm|9819/3|Leukemia__B_Cell
C019|Root_Of_Tongue|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C019|Root_Of_Tongue|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C019|Root_Of_Tongue|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C019|Root_Of_Tongue|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C019|Root_Of_Tongue|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C019|Root_Of_Tongue|997|Neoplasm|9971/3|Polymorphic_PTLD
C019|Root_Of_Tongue|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C020-C024,C028-C029|Root_Of_Tongue|800|Neoplasm|8000/3|Malignant_Neoplasm
C020-C024,C028-C029|Root_Of_Tongue|800|Neoplasm|8001/3|Malignant_Cell
C020-C024,C028-C029|Root_Of_Tongue|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C020-C024,C028-C029|Root_Of_Tongue|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C020-C024,C028-C029|Root_Of_Tongue|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C020-C024,C028-C029|Root_Of_Tongue|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C020-C024,C028-C029|Root_Of_Tongue|801|Carcinoma|8010/2|In_Situ_Cancer
C020-C024,C028-C029|Root_Of_Tongue|801|Carcinoma|8010/3|Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|801|Carcinoma|8011/3|Malignant_Epithelioma
C020-C024,C028-C029|Root_Of_Tongue|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C020-C024,C028-C029|Root_Of_Tongue|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C020-C024,C028-C029|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C020-C024,C028-C029|Root_Of_Tongue|814|Adenocarcinoma|8140/3|Adenocarcinoma
C020-C024,C028-C029|Root_Of_Tongue|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C020-C024,C028-C029|Root_Of_Tongue|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C020-C024,C028-C029|Root_Of_Tongue|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C020-C024,C028-C029|Root_Of_Tongue|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C020-C024,C028-C029|Root_Of_Tongue|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C020-C024,C028-C029|Root_Of_Tongue|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C020-C024,C028-C029|Root_Of_Tongue|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C020-C024,C028-C029|Root_Of_Tongue|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C020-C024,C028-C029|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C020-C024,C028-C029|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C020-C024,C028-C029|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C020-C024,C028-C029|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C020-C024,C028-C029|Root_Of_Tongue|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C020-C024,C028-C029|Root_Of_Tongue|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C020-C024,C028-C029|Root_Of_Tongue|872|Melanoma|8720/3|Melanoma
C020-C024,C028-C029|Root_Of_Tongue|872|Melanoma|8721/3|Nodular_Melanoma
C020-C024,C028-C029|Root_Of_Tongue|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C020-C024,C028-C029|Root_Of_Tongue|872|Melanoma|8723/3|Regressing_Melanoma
C020-C024,C028-C029|Root_Of_Tongue|882|Sarcoma|8825/3|Sarcoma
C020-C024,C028-C029|Root_Of_Tongue|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C020-C024,C028-C029|Root_Of_Tongue|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C020-C024,C028-C029|Root_Of_Tongue|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C020-C024,C028-C029|Root_Of_Tongue|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C020-C024,C028-C029|Root_Of_Tongue|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C020-C024,C028-C029|Root_Of_Tongue|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C020-C024,C028-C029|Root_Of_Tongue|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C020-C024,C028-C029|Root_Of_Tongue|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C020-C024,C028-C029|Root_Of_Tongue|959|Lymphoma|9590/3|Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C020-C024,C028-C029|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C020-C024,C028-C029|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C020-C024,C028-C029|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C020-C024,C028-C029|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C020-C024,C028-C029|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C020-C024,C028-C029|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C020-C024,C028-C029|Root_Of_Tongue|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C020-C024,C028-C029|Root_Of_Tongue|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C020-C024,C028-C029|Root_Of_Tongue|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C020-C024,C028-C029|Root_Of_Tongue|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C020-C024,C028-C029|Root_Of_Tongue|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C020-C024,C028-C029|Root_Of_Tongue|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C020-C024,C028-C029|Root_Of_Tongue|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|973|Plasmacytoma|9731/3|Plasmacytoma
C020-C024,C028-C029|Root_Of_Tongue|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C020-C024,C028-C029|Root_Of_Tongue|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C020-C024,C028-C029|Root_Of_Tongue|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C020-C024,C028-C029|Root_Of_Tongue|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C020-C024,C028-C029|Root_Of_Tongue|975|Neoplasm|9750/3|Malignant_Histiocytosis
C020-C024,C028-C029|Root_Of_Tongue|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C020-C024,C028-C029|Root_Of_Tongue|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C020-C024,C028-C029|Root_Of_Tongue|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C020-C024,C028-C029|Root_Of_Tongue|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C020-C024,C028-C029|Root_Of_Tongue|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C020-C024,C028-C029|Root_Of_Tongue|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C020-C024,C028-C029|Root_Of_Tongue|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C020-C024,C028-C029|Root_Of_Tongue|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9812/3|Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9813/3|Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9814/3|Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9816/3|Hypodiploid_ALL
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9817/3|Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9818/3|Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|981|Neoplasm|9819/3|Leukemia__B_Cell
C020-C024,C028-C029|Root_Of_Tongue|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C020-C024,C028-C029|Root_Of_Tongue|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C020-C024,C028-C029|Root_Of_Tongue|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C020-C024,C028-C029|Root_Of_Tongue|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C020-C024,C028-C029|Root_Of_Tongue|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C020-C024,C028-C029|Root_Of_Tongue|997|Neoplasm|9971/3|Polymorphic_PTLD
C020-C024,C028-C029|Root_Of_Tongue|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|800|Neoplasm|8000/3|Malignant_Neoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|800|Neoplasm|8001/3|Malignant_Cell
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|801|Carcinoma|8010/2|In_Situ_Cancer
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|801|Carcinoma|8010/3|Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|801|Carcinoma|8011/3|Malignant_Epithelioma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|814|Adenocarcinoma|8140/3|Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|872|Melanoma|8720/3|Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|872|Melanoma|8721/3|Nodular_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|872|Melanoma|8723/3|Regressing_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|874|Nevus|8745/3|Desmoplastic_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|882|Sarcoma|8825/3|Sarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|898|Carcinosarcoma|8980/3|Carcinosarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|959|Lymphoma|9590/3|Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|973|Plasmacytoma|9731/3|Plasmacytoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|975|Neoplasm|9750/3|Malignant_Histiocytosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9812/3|Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9813/3|Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9814/3|Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9816/3|Hypodiploid_ALL
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9817/3|Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9818/3|Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|981|Neoplasm|9819/3|Leukemia__B_Cell
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|997|Neoplasm|9971/3|Polymorphic_PTLD
C030-C031,C039-C041,C048-C052,C058-C062,C068-C069|Sublingual_Region|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C079-C081,C088-C089|Salivary_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C079-C081,C088-C089|Salivary_Gland|800|Neoplasm|8001/3|Malignant_Cell
C079-C081,C088-C089|Salivary_Gland|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C079-C081,C088-C089|Salivary_Gland|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C079-C081,C088-C089|Salivary_Gland|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C079-C081,C088-C089|Salivary_Gland|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C079-C081,C088-C089|Salivary_Gland|801|Carcinoma|8010/2|In_Situ_Cancer
C079-C081,C088-C089|Salivary_Gland|801|Carcinoma|8010/3|Carcinoma
C079-C081,C088-C089|Salivary_Gland|801|Carcinoma|8011/3|Malignant_Epithelioma
C079-C081,C088-C089|Salivary_Gland|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C079-C081,C088-C089|Salivary_Gland|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C079-C081,C088-C089|Salivary_Gland|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C079-C081,C088-C089|Salivary_Gland|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C079-C081,C088-C089|Salivary_Gland|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C079-C081,C088-C089|Salivary_Gland|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C079-C081,C088-C089|Salivary_Gland|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C079-C081,C088-C089|Salivary_Gland|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C079-C081,C088-C089|Salivary_Gland|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C079-C081,C088-C089|Salivary_Gland|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C079-C081,C088-C089|Salivary_Gland|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C079-C081,C088-C089|Salivary_Gland|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C079-C081,C088-C089|Salivary_Gland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C079-C081,C088-C089|Salivary_Gland|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C079-C081,C088-C089|Salivary_Gland|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C079-C081,C088-C089|Salivary_Gland|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C079-C081,C088-C089|Salivary_Gland|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C079-C081,C088-C089|Salivary_Gland|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C079-C081,C088-C089|Salivary_Gland|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C079-C081,C088-C089|Salivary_Gland|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C079-C081,C088-C089|Salivary_Gland|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C079-C081,C088-C089|Salivary_Gland|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C079-C081,C088-C089|Salivary_Gland|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C079-C081,C088-C089|Salivary_Gland|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C079-C081,C088-C089|Salivary_Gland|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C079-C081,C088-C089|Salivary_Gland|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C079-C081,C088-C089|Salivary_Gland|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|850|Ductal_Carcinoma|8500/3|Invasive_Carcinoma
C079-C081,C088-C089|Salivary_Gland|850|Ductal_Carcinoma|8502/3|Secretory_Breast_Carcinoma
C079-C081,C088-C089|Salivary_Gland|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C079-C081,C088-C089|Salivary_Gland|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C079-C081,C088-C089|Salivary_Gland|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C079-C081,C088-C089|Salivary_Gland|856|Adenosquamous_Carcinoma|8561/3|Malignant_Neoplasm
C079-C081,C088-C089|Salivary_Gland|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C079-C081,C088-C089|Salivary_Gland|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C079-C081,C088-C089|Salivary_Gland|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C079-C081,C088-C089|Salivary_Gland|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C079-C081,C088-C089|Salivary_Gland|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C079-C081,C088-C089|Salivary_Gland|880|Sarcoma|8800/3|Sarcoma
C079-C081,C088-C089|Salivary_Gland|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C079-C081,C088-C089|Salivary_Gland|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C079-C081,C088-C089|Salivary_Gland|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C079-C081,C088-C089|Salivary_Gland|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C079-C081,C088-C089|Salivary_Gland|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C079-C081,C088-C089|Salivary_Gland|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C079-C081,C088-C089|Salivary_Gland|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C079-C081,C088-C089|Salivary_Gland|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C079-C081,C088-C089|Salivary_Gland|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C079-C081,C088-C089|Salivary_Gland|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C079-C081,C088-C089|Salivary_Gland|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C079-C081,C088-C089|Salivary_Gland|882|Sarcoma|8825/3|Sarcoma
C079-C081,C088-C089|Salivary_Gland|884|Myxosarcoma|8840/3|Myxosarcoma
C079-C081,C088-C089|Salivary_Gland|885|Liposarcoma|8850/3|Liposarcoma
C079-C081,C088-C089|Salivary_Gland|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C079-C081,C088-C089|Salivary_Gland|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C079-C081,C088-C089|Salivary_Gland|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C079-C081,C088-C089|Salivary_Gland|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C079-C081,C088-C089|Salivary_Gland|885|Liposarcoma|8855/3|Liposarcoma
C079-C081,C088-C089|Salivary_Gland|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C079-C081,C088-C089|Salivary_Gland|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C079-C081,C088-C089|Salivary_Gland|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C079-C081,C088-C089|Salivary_Gland|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C079-C081,C088-C089|Salivary_Gland|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C079-C081,C088-C089|Salivary_Gland|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C079-C081,C088-C089|Salivary_Gland|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C079-C081,C088-C089|Salivary_Gland|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C079-C081,C088-C089|Salivary_Gland|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C079-C081,C088-C089|Salivary_Gland|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C079-C081,C088-C089|Salivary_Gland|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C079-C081,C088-C089|Salivary_Gland|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C079-C081,C088-C089|Salivary_Gland|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C079-C081,C088-C089|Salivary_Gland|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C079-C081,C088-C089|Salivary_Gland|898|Carcinosarcoma|8980/3|Carcinosarcoma
C079-C081,C088-C089|Salivary_Gland|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C079-C081,C088-C089|Salivary_Gland|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C079-C081,C088-C089|Salivary_Gland|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C079-C081,C088-C089|Salivary_Gland|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C079-C081,C088-C089|Salivary_Gland|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C079-C081,C088-C089|Salivary_Gland|959|Lymphoma|9590/3|Lymphoma
C079-C081,C088-C089|Salivary_Gland|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C079-C081,C088-C089|Salivary_Gland|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C079-C081,C088-C089|Salivary_Gland|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C079-C081,C088-C089|Salivary_Gland|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C079-C081,C088-C089|Salivary_Gland|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C079-C081,C088-C089|Salivary_Gland|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C079-C081,C088-C089|Salivary_Gland|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C079-C081,C088-C089|Salivary_Gland|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C079-C081,C088-C089|Salivary_Gland|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C079-C081,C088-C089|Salivary_Gland|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C079-C081,C088-C089|Salivary_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C079-C081,C088-C089|Salivary_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C079-C081,C088-C089|Salivary_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C079-C081,C088-C089|Salivary_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C079-C081,C088-C089|Salivary_Gland|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C079-C081,C088-C089|Salivary_Gland|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C079-C081,C088-C089|Salivary_Gland|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C079-C081,C088-C089|Salivary_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C079-C081,C088-C089|Salivary_Gland|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C079-C081,C088-C089|Salivary_Gland|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C079-C081,C088-C089|Salivary_Gland|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C079-C081,C088-C089|Salivary_Gland|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C079-C081,C088-C089|Salivary_Gland|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C079-C081,C088-C089|Salivary_Gland|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C079-C081,C088-C089|Salivary_Gland|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C079-C081,C088-C089|Salivary_Gland|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C079-C081,C088-C089|Salivary_Gland|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C079-C081,C088-C089|Salivary_Gland|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C079-C081,C088-C089|Salivary_Gland|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C079-C081,C088-C089|Salivary_Gland|973|Plasmacytoma|9731/3|Plasmacytoma
C079-C081,C088-C089|Salivary_Gland|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C079-C081,C088-C089|Salivary_Gland|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C079-C081,C088-C089|Salivary_Gland|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C079-C081,C088-C089|Salivary_Gland|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C079-C081,C088-C089|Salivary_Gland|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C079-C081,C088-C089|Salivary_Gland|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C079-C081,C088-C089|Salivary_Gland|975|Neoplasm|9750/3|Malignant_Histiocytosis
C079-C081,C088-C089|Salivary_Gland|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C079-C081,C088-C089|Salivary_Gland|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C079-C081,C088-C089|Salivary_Gland|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C079-C081,C088-C089|Salivary_Gland|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C079-C081,C088-C089|Salivary_Gland|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C079-C081,C088-C089|Salivary_Gland|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C079-C081,C088-C089|Salivary_Gland|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C079-C081,C088-C089|Salivary_Gland|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9812/3|Lymphoma
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9813/3|Lymphoma
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9814/3|Lymphoma
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9816/3|Hypodiploid_ALL
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9817/3|Lymphoma
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9818/3|Lymphoma
C079-C081,C088-C089|Salivary_Gland|981|Neoplasm|9819/3|Leukemia__B_Cell
C079-C081,C088-C089|Salivary_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C079-C081,C088-C089|Salivary_Gland|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C079-C081,C088-C089|Salivary_Gland|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C079-C081,C088-C089|Salivary_Gland|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C079-C081,C088-C089|Salivary_Gland|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C079-C081,C088-C089|Salivary_Gland|997|Neoplasm|9971/3|Polymorphic_PTLD
C079-C081,C088-C089|Salivary_Gland|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C090-C091,C098-C104,C108-C109|Pharynx|800|Neoplasm|8000/3|Malignant_Neoplasm
C090-C091,C098-C104,C108-C109|Pharynx|800|Neoplasm|8001/3|Malignant_Cell
C090-C091,C098-C104,C108-C109|Pharynx|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C090-C091,C098-C104,C108-C109|Pharynx|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C090-C091,C098-C104,C108-C109|Pharynx|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C090-C091,C098-C104,C108-C109|Pharynx|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8010/2|In_Situ_Cancer
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8010/3|Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8011/3|Malignant_Epithelioma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C090-C091,C098-C104,C108-C109|Pharynx|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C090-C091,C098-C104,C108-C109|Pharynx|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|Lymphoepithelial_Carcinoma|8085/3|Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|808|Lymphoepithelial_Carcinoma|8086/3|Squamous_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C090-C091,C098-C104,C108-C109|Pharynx|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C090-C091,C098-C104,C108-C109|Pharynx|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C090-C091,C098-C104,C108-C109|Pharynx|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C090-C091,C098-C104,C108-C109|Pharynx|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C090-C091,C098-C104,C108-C109|Pharynx|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C090-C091,C098-C104,C108-C109|Pharynx|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C090-C091,C098-C104,C108-C109|Pharynx|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C090-C091,C098-C104,C108-C109|Pharynx|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8720/3|Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8721/3|Nodular_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|872|Melanoma|8723/3|Regressing_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C090-C091,C098-C104,C108-C109|Pharynx|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|874|Nevus|8745/3|Desmoplastic_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|876|Nevus|8761/3|Giant_Congenital_Nevus
C090-C091,C098-C104,C108-C109|Pharynx|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8800/3|Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8850/3|Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8855/3|Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C090-C091,C098-C104,C108-C109|Pharynx|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C090-C091,C098-C104,C108-C109|Pharynx|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C090-C091,C098-C104,C108-C109|Pharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C090-C091,C098-C104,C108-C109|Pharynx|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C090-C091,C098-C104,C108-C109|Pharynx|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C090-C091,C098-C104,C108-C109|Pharynx|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|959|Lymphoma|9590/3|Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C090-C091,C098-C104,C108-C109|Pharynx|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C090-C091,C098-C104,C108-C109|Pharynx|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C090-C091,C098-C104,C108-C109|Pharynx|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C090-C091,C098-C104,C108-C109|Pharynx|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C090-C091,C098-C104,C108-C109|Pharynx|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C090-C091,C098-C104,C108-C109|Pharynx|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C090-C091,C098-C104,C108-C109|Pharynx|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C090-C091,C098-C104,C108-C109|Pharynx|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C090-C091,C098-C104,C108-C109|Pharynx|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C090-C091,C098-C104,C108-C109|Pharynx|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C090-C091,C098-C104,C108-C109|Pharynx|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C090-C091,C098-C104,C108-C109|Pharynx|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C090-C091,C098-C104,C108-C109|Pharynx|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C090-C091,C098-C104,C108-C109|Pharynx|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C090-C091,C098-C104,C108-C109|Pharynx|975|Neoplasm|9750/3|Malignant_Histiocytosis
C090-C091,C098-C104,C108-C109|Pharynx|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C090-C091,C098-C104,C108-C109|Pharynx|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C090-C091,C098-C104,C108-C109|Pharynx|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C090-C091,C098-C104,C108-C109|Pharynx|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C090-C091,C098-C104,C108-C109|Pharynx|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9812/3|Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9813/3|Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9814/3|Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9816/3|Hypodiploid_ALL
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9817/3|Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9818/3|Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|981|Neoplasm|9819/3|Leukemia__B_Cell
C090-C091,C098-C104,C108-C109|Pharynx|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C090-C091,C098-C104,C108-C109|Pharynx|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C090-C091,C098-C104,C108-C109|Pharynx|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C090-C091,C098-C104,C108-C109|Pharynx|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C090-C091,C098-C104,C108-C109|Pharynx|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C090-C091,C098-C104,C108-C109|Pharynx|997|Neoplasm|9971/3|Polymorphic_PTLD
C090-C091,C098-C104,C108-C109|Pharynx|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C110,C112-C113,C118-C119|Nasopharynx|800|Neoplasm|8000/3|Malignant_Neoplasm
C110,C112-C113,C118-C119|Nasopharynx|800|Neoplasm|8001/3|Malignant_Cell
C110,C112-C113,C118-C119|Nasopharynx|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C110,C112-C113,C118-C119|Nasopharynx|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C110,C112-C113,C118-C119|Nasopharynx|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C110,C112-C113,C118-C119|Nasopharynx|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8010/2|In_Situ_Cancer
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8010/3|Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8011/3|Malignant_Epithelioma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C110,C112-C113,C118-C119|Nasopharynx|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C110,C112-C113,C118-C119|Nasopharynx|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C110,C112-C113,C118-C119|Nasopharynx|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C110,C112-C113,C118-C119|Nasopharynx|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C110,C112-C113,C118-C119|Nasopharynx|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C110,C112-C113,C118-C119|Nasopharynx|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C110,C112-C113,C118-C119|Nasopharynx|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C110,C112-C113,C118-C119|Nasopharynx|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C110,C112-C113,C118-C119|Nasopharynx|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C110,C112-C113,C118-C119|Nasopharynx|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8720/3|Melanoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8721/3|Nodular_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|872|Melanoma|8723/3|Regressing_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C110,C112-C113,C118-C119|Nasopharynx|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|874|Nevus|8745/3|Desmoplastic_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8800/3|Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C110,C112-C113,C118-C119|Nasopharynx|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C110,C112-C113,C118-C119|Nasopharynx|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C110,C112-C113,C118-C119|Nasopharynx|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C110,C112-C113,C118-C119|Nasopharynx|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C110,C112-C113,C118-C119|Nasopharynx|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C110,C112-C113,C118-C119|Nasopharynx|882|Sarcoma|8825/3|Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C110,C112-C113,C118-C119|Nasopharynx|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C110,C112-C113,C118-C119|Nasopharynx|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C110,C112-C113,C118-C119|Nasopharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C110,C112-C113,C118-C119|Nasopharynx|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C110,C112-C113,C118-C119|Nasopharynx|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C110,C112-C113,C118-C119|Nasopharynx|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C110,C112-C113,C118-C119|Nasopharynx|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C110,C112-C113,C118-C119|Nasopharynx|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C110,C112-C113,C118-C119|Nasopharynx|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|937|Chordoma|9370/3|Chordoma
C110,C112-C113,C118-C119|Nasopharynx|937|Chordoma|9371/3|Chondroid_Chordoma
C110,C112-C113,C118-C119|Nasopharynx|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C110,C112-C113,C118-C119|Nasopharynx|959|Lymphoma|9590/3|Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C110,C112-C113,C118-C119|Nasopharynx|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C110,C112-C113,C118-C119|Nasopharynx|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C110,C112-C113,C118-C119|Nasopharynx|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C110,C112-C113,C118-C119|Nasopharynx|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C110,C112-C113,C118-C119|Nasopharynx|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C110,C112-C113,C118-C119|Nasopharynx|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C110,C112-C113,C118-C119|Nasopharynx|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C110,C112-C113,C118-C119|Nasopharynx|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C110,C112-C113,C118-C119|Nasopharynx|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C110,C112-C113,C118-C119|Nasopharynx|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C110,C112-C113,C118-C119|Nasopharynx|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C110,C112-C113,C118-C119|Nasopharynx|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C110,C112-C113,C118-C119|Nasopharynx|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C110,C112-C113,C118-C119|Nasopharynx|975|Neoplasm|9750/3|Malignant_Histiocytosis
C110,C112-C113,C118-C119|Nasopharynx|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C110,C112-C113,C118-C119|Nasopharynx|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C110,C112-C113,C118-C119|Nasopharynx|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C110,C112-C113,C118-C119|Nasopharynx|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C110,C112-C113,C118-C119|Nasopharynx|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9812/3|Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9813/3|Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9814/3|Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9816/3|Hypodiploid_ALL
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9817/3|Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9818/3|Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|981|Neoplasm|9819/3|Leukemia__B_Cell
C110,C112-C113,C118-C119|Nasopharynx|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C110,C112-C113,C118-C119|Nasopharynx|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C110,C112-C113,C118-C119|Nasopharynx|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C110,C112-C113,C118-C119|Nasopharynx|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C110,C112-C113,C118-C119|Nasopharynx|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C110,C112-C113,C118-C119|Nasopharynx|997|Neoplasm|9971/3|Polymorphic_PTLD
C110,C112-C113,C118-C119|Nasopharynx|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C111|Posterior_Wall_Of_The_Nasopharynx|800|Neoplasm|8000/3|Malignant_Neoplasm
C111|Posterior_Wall_Of_The_Nasopharynx|800|Neoplasm|8001/3|Malignant_Cell
C111|Posterior_Wall_Of_The_Nasopharynx|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C111|Posterior_Wall_Of_The_Nasopharynx|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C111|Posterior_Wall_Of_The_Nasopharynx|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C111|Posterior_Wall_Of_The_Nasopharynx|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C111|Posterior_Wall_Of_The_Nasopharynx|801|Carcinoma|8010/2|In_Situ_Cancer
C111|Posterior_Wall_Of_The_Nasopharynx|801|Carcinoma|8010/3|Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|801|Carcinoma|8011/3|Malignant_Epithelioma
C111|Posterior_Wall_Of_The_Nasopharynx|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C111|Posterior_Wall_Of_The_Nasopharynx|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C111|Posterior_Wall_Of_The_Nasopharynx|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C111|Posterior_Wall_Of_The_Nasopharynx|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|808|Lymphoepithelial_Carcinoma|8085/3|Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|808|Lymphoepithelial_Carcinoma|8086/3|Squamous_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C111|Posterior_Wall_Of_The_Nasopharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C111|Posterior_Wall_Of_The_Nasopharynx|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C111|Posterior_Wall_Of_The_Nasopharynx|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C111|Posterior_Wall_Of_The_Nasopharynx|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C111|Posterior_Wall_Of_The_Nasopharynx|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C111|Posterior_Wall_Of_The_Nasopharynx|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C111|Posterior_Wall_Of_The_Nasopharynx|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C111|Posterior_Wall_Of_The_Nasopharynx|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|872|Melanoma|8720/3|Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|872|Melanoma|8721/3|Nodular_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|872|Melanoma|8723/3|Regressing_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C111|Posterior_Wall_Of_The_Nasopharynx|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|874|Nevus|8745/3|Desmoplastic_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C111|Posterior_Wall_Of_The_Nasopharynx|880|Sarcoma|8800/3|Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C111|Posterior_Wall_Of_The_Nasopharynx|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C111|Posterior_Wall_Of_The_Nasopharynx|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C111|Posterior_Wall_Of_The_Nasopharynx|882|Sarcoma|8825/3|Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C111|Posterior_Wall_Of_The_Nasopharynx|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C111|Posterior_Wall_Of_The_Nasopharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C111|Posterior_Wall_Of_The_Nasopharynx|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C111|Posterior_Wall_Of_The_Nasopharynx|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C111|Posterior_Wall_Of_The_Nasopharynx|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C111|Posterior_Wall_Of_The_Nasopharynx|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C111|Posterior_Wall_Of_The_Nasopharynx|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|937|Chordoma|9370/3|Chordoma
C111|Posterior_Wall_Of_The_Nasopharynx|937|Chordoma|9371/3|Chondroid_Chordoma
C111|Posterior_Wall_Of_The_Nasopharynx|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C111|Posterior_Wall_Of_The_Nasopharynx|959|Lymphoma|9590/3|Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C111|Posterior_Wall_Of_The_Nasopharynx|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C111|Posterior_Wall_Of_The_Nasopharynx|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C111|Posterior_Wall_Of_The_Nasopharynx|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C111|Posterior_Wall_Of_The_Nasopharynx|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C111|Posterior_Wall_Of_The_Nasopharynx|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C111|Posterior_Wall_Of_The_Nasopharynx|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C111|Posterior_Wall_Of_The_Nasopharynx|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C111|Posterior_Wall_Of_The_Nasopharynx|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C111|Posterior_Wall_Of_The_Nasopharynx|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C111|Posterior_Wall_Of_The_Nasopharynx|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C111|Posterior_Wall_Of_The_Nasopharynx|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C111|Posterior_Wall_Of_The_Nasopharynx|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C111|Posterior_Wall_Of_The_Nasopharynx|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C111|Posterior_Wall_Of_The_Nasopharynx|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C111|Posterior_Wall_Of_The_Nasopharynx|975|Neoplasm|9750/3|Malignant_Histiocytosis
C111|Posterior_Wall_Of_The_Nasopharynx|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C111|Posterior_Wall_Of_The_Nasopharynx|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C111|Posterior_Wall_Of_The_Nasopharynx|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C111|Posterior_Wall_Of_The_Nasopharynx|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C111|Posterior_Wall_Of_The_Nasopharynx|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|981|Neoplasm|9812/3|Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|981|Neoplasm|9813/3|Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|981|Neoplasm|9814/3|Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|981|Neoplasm|9816/3|Hypodiploid_ALL
C111|Posterior_Wall_Of_The_Nasopharynx|981|Neoplasm|9817/3|Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|981|Neoplasm|9818/3|Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C111|Posterior_Wall_Of_The_Nasopharynx|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C111|Posterior_Wall_Of_The_Nasopharynx|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C111|Posterior_Wall_Of_The_Nasopharynx|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C111|Posterior_Wall_Of_The_Nasopharynx|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C111|Posterior_Wall_Of_The_Nasopharynx|997|Neoplasm|9971/3|Polymorphic_PTLD
C111|Posterior_Wall_Of_The_Nasopharynx|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C129-C132,C138-C139|Hypopharynx|800|Neoplasm|8000/3|Malignant_Neoplasm
C129-C132,C138-C139|Hypopharynx|800|Neoplasm|8001/3|Malignant_Cell
C129-C132,C138-C139|Hypopharynx|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C129-C132,C138-C139|Hypopharynx|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C129-C132,C138-C139|Hypopharynx|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C129-C132,C138-C139|Hypopharynx|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8010/2|In_Situ_Cancer
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8010/3|Carcinoma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8011/3|Malignant_Epithelioma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C129-C132,C138-C139|Hypopharynx|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C129-C132,C138-C139|Hypopharynx|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C129-C132,C138-C139|Hypopharynx|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C129-C132,C138-C139|Hypopharynx|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C129-C132,C138-C139|Hypopharynx|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C129-C132,C138-C139|Hypopharynx|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C129-C132,C138-C139|Hypopharynx|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C129-C132,C138-C139|Hypopharynx|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C129-C132,C138-C139|Hypopharynx|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C129-C132,C138-C139|Hypopharynx|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C129-C132,C138-C139|Hypopharynx|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C129-C132,C138-C139|Hypopharynx|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C129-C132,C138-C139|Hypopharynx|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C129-C132,C138-C139|Hypopharynx|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C129-C132,C138-C139|Hypopharynx|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C129-C132,C138-C139|Hypopharynx|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C129-C132,C138-C139|Hypopharynx|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C129-C132,C138-C139|Hypopharynx|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C129-C132,C138-C139|Hypopharynx|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C129-C132,C138-C139|Hypopharynx|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C129-C132,C138-C139|Hypopharynx|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C129-C132,C138-C139|Hypopharynx|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C129-C132,C138-C139|Hypopharynx|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C129-C132,C138-C139|Hypopharynx|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C129-C132,C138-C139|Hypopharynx|882|Sarcoma|8825/3|Sarcoma
C129-C132,C138-C139|Hypopharynx|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C129-C132,C138-C139|Hypopharynx|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C129-C132,C138-C139|Hypopharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C129-C132,C138-C139|Hypopharynx|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C129-C132,C138-C139|Hypopharynx|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C129-C132,C138-C139|Hypopharynx|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C129-C132,C138-C139|Hypopharynx|959|Lymphoma|9590/3|Lymphoma
C129-C132,C138-C139|Hypopharynx|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C129-C132,C138-C139|Hypopharynx|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C129-C132,C138-C139|Hypopharynx|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C129-C132,C138-C139|Hypopharynx|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C129-C132,C138-C139|Hypopharynx|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C129-C132,C138-C139|Hypopharynx|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C129-C132,C138-C139|Hypopharynx|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C129-C132,C138-C139|Hypopharynx|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C129-C132,C138-C139|Hypopharynx|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C129-C132,C138-C139|Hypopharynx|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C129-C132,C138-C139|Hypopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C129-C132,C138-C139|Hypopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C129-C132,C138-C139|Hypopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C129-C132,C138-C139|Hypopharynx|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C129-C132,C138-C139|Hypopharynx|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C129-C132,C138-C139|Hypopharynx|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C129-C132,C138-C139|Hypopharynx|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C129-C132,C138-C139|Hypopharynx|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C129-C132,C138-C139|Hypopharynx|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C129-C132,C138-C139|Hypopharynx|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C129-C132,C138-C139|Hypopharynx|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C129-C132,C138-C139|Hypopharynx|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C129-C132,C138-C139|Hypopharynx|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C129-C132,C138-C139|Hypopharynx|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C129-C132,C138-C139|Hypopharynx|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C129-C132,C138-C139|Hypopharynx|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C129-C132,C138-C139|Hypopharynx|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C129-C132,C138-C139|Hypopharynx|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C129-C132,C138-C139|Hypopharynx|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C129-C132,C138-C139|Hypopharynx|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C129-C132,C138-C139|Hypopharynx|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C129-C132,C138-C139|Hypopharynx|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C129-C132,C138-C139|Hypopharynx|975|Neoplasm|9750/3|Malignant_Histiocytosis
C129-C132,C138-C139|Hypopharynx|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C129-C132,C138-C139|Hypopharynx|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C129-C132,C138-C139|Hypopharynx|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C129-C132,C138-C139|Hypopharynx|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C129-C132,C138-C139|Hypopharynx|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C129-C132,C138-C139|Hypopharynx|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C129-C132,C138-C139|Hypopharynx|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C129-C132,C138-C139|Hypopharynx|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9812/3|Lymphoma
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9813/3|Lymphoma
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9814/3|Lymphoma
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9816/3|Hypodiploid_ALL
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9817/3|Lymphoma
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9818/3|Lymphoma
C129-C132,C138-C139|Hypopharynx|981|Neoplasm|9819/3|Leukemia__B_Cell
C129-C132,C138-C139|Hypopharynx|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C129-C132,C138-C139|Hypopharynx|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C129-C132,C138-C139|Hypopharynx|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C129-C132,C138-C139|Hypopharynx|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C129-C132,C138-C139|Hypopharynx|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C129-C132,C138-C139|Hypopharynx|997|Neoplasm|9971/3|Polymorphic_PTLD
C129-C132,C138-C139|Hypopharynx|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C140,C142,C148|Pharynx|800|Neoplasm|8000/3|Malignant_Neoplasm
C140,C142,C148|Pharynx|800|Neoplasm|8001/3|Malignant_Cell
C140,C142,C148|Pharynx|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C140,C142,C148|Pharynx|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C140,C142,C148|Pharynx|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C140,C142,C148|Pharynx|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C140,C142,C148|Pharynx|801|Carcinoma|8010/2|In_Situ_Cancer
C140,C142,C148|Pharynx|801|Carcinoma|8010/3|Carcinoma
C140,C142,C148|Pharynx|801|Carcinoma|8011/3|Malignant_Epithelioma
C140,C142,C148|Pharynx|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C140,C142,C148|Pharynx|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C140,C142,C148|Pharynx|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C140,C142,C148|Pharynx|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C140,C142,C148|Pharynx|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C140,C142,C148|Pharynx|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C140,C142,C148|Pharynx|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C140,C142,C148|Pharynx|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C140,C142,C148|Pharynx|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C140,C142,C148|Pharynx|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C140,C142,C148|Pharynx|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C140,C142,C148|Pharynx|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C140,C142,C148|Pharynx|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C140,C142,C148|Pharynx|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C140,C142,C148|Pharynx|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C140,C142,C148|Pharynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C140,C142,C148|Pharynx|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C140,C142,C148|Pharynx|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C140,C142,C148|Pharynx|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C140,C142,C148|Pharynx|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C140,C142,C148|Pharynx|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C140,C142,C148|Pharynx|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C140,C142,C148|Pharynx|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C140,C142,C148|Pharynx|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C140,C142,C148|Pharynx|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C140,C142,C148|Pharynx|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C140,C142,C148|Pharynx|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C140,C142,C148|Pharynx|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C140,C142,C148|Pharynx|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C140,C142,C148|Pharynx|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C140,C142,C148|Pharynx|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C140,C142,C148|Pharynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C140,C142,C148|Pharynx|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C140,C142,C148|Pharynx|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C140,C142,C148|Pharynx|937|Chordoma|9370/3|Chordoma
C140,C142,C148|Pharynx|937|Chordoma|9371/3|Chondroid_Chordoma
C140,C142,C148|Pharynx|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C140,C142,C148|Pharynx|959|Lymphoma|9590/3|Lymphoma
C140,C142,C148|Pharynx|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C140,C142,C148|Pharynx|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C140,C142,C148|Pharynx|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C140,C142,C148|Pharynx|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C140,C142,C148|Pharynx|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C140,C142,C148|Pharynx|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C140,C142,C148|Pharynx|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C140,C142,C148|Pharynx|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C140,C142,C148|Pharynx|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C140,C142,C148|Pharynx|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C140,C142,C148|Pharynx|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C140,C142,C148|Pharynx|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C140,C142,C148|Pharynx|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C140,C142,C148|Pharynx|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C140,C142,C148|Pharynx|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C140,C142,C148|Pharynx|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C140,C142,C148|Pharynx|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C140,C142,C148|Pharynx|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C140,C142,C148|Pharynx|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C140,C142,C148|Pharynx|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C140,C142,C148|Pharynx|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C140,C142,C148|Pharynx|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C140,C142,C148|Pharynx|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C140,C142,C148|Pharynx|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C140,C142,C148|Pharynx|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C140,C142,C148|Pharynx|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C140,C142,C148|Pharynx|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C140,C142,C148|Pharynx|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C140,C142,C148|Pharynx|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9731/3|Plasmacytoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C140,C142,C148|Pharynx|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C140,C142,C148|Pharynx|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C140,C142,C148|Pharynx|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C140,C142,C148|Pharynx|975|Neoplasm|9750/3|Malignant_Histiocytosis
C140,C142,C148|Pharynx|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C140,C142,C148|Pharynx|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C140,C142,C148|Pharynx|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C140,C142,C148|Pharynx|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C140,C142,C148|Pharynx|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C140,C142,C148|Pharynx|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C140,C142,C148|Pharynx|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C140,C142,C148|Pharynx|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C140,C142,C148|Pharynx|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C140,C142,C148|Pharynx|981|Neoplasm|9812/3|Lymphoma
C140,C142,C148|Pharynx|981|Neoplasm|9813/3|Lymphoma
C140,C142,C148|Pharynx|981|Neoplasm|9814/3|Lymphoma
C140,C142,C148|Pharynx|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C140,C142,C148|Pharynx|981|Neoplasm|9816/3|Hypodiploid_ALL
C140,C142,C148|Pharynx|981|Neoplasm|9817/3|Lymphoma
C140,C142,C148|Pharynx|981|Neoplasm|9818/3|Lymphoma
C140,C142,C148|Pharynx|981|Neoplasm|9819/3|Leukemia__B_Cell
C140,C142,C148|Pharynx|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C140,C142,C148|Pharynx|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C140,C142,C148|Pharynx|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C140,C142,C148|Pharynx|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C140,C142,C148|Pharynx|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C140,C142,C148|Pharynx|997|Neoplasm|9971/3|Polymorphic_PTLD
C140,C142,C148|Pharynx|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C150-C155,C158-C159|Esophagus|800|Neoplasm|8000/3|Malignant_Neoplasm
C150-C155,C158-C159|Esophagus|800|Neoplasm|8001/3|Malignant_Cell
C150-C155,C158-C159|Esophagus|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C150-C155,C158-C159|Esophagus|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C150-C155,C158-C159|Esophagus|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C150-C155,C158-C159|Esophagus|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C150-C155,C158-C159|Esophagus|801|Carcinoma|8010/2|In_Situ_Cancer
C150-C155,C158-C159|Esophagus|801|Carcinoma|8010/3|Carcinoma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8011/3|Malignant_Epithelioma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C150-C155,C158-C159|Esophagus|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C150-C155,C158-C159|Esophagus|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C150-C155,C158-C159|Esophagus|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C150-C155,C158-C159|Esophagus|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C150-C155,C158-C159|Esophagus|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C150-C155,C158-C159|Esophagus|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C150-C155,C158-C159|Esophagus|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C150-C155,C158-C159|Esophagus|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C150-C155,C158-C159|Esophagus|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C150-C155,C158-C159|Esophagus|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C150-C155,C158-C159|Esophagus|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8145/3|Diffuse_Type_Adenocarcinoma
C150-C155,C158-C159|Esophagus|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C150-C155,C158-C159|Esophagus|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C150-C155,C158-C159|Esophagus|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C150-C155,C158-C159|Esophagus|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C150-C155,C158-C159|Esophagus|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C150-C155,C158-C159|Esophagus|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C150-C155,C158-C159|Esophagus|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C150-C155,C158-C159|Esophagus|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C150-C155,C158-C159|Esophagus|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C150-C155,C158-C159|Esophagus|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C150-C155,C158-C159|Esophagus|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C150-C155,C158-C159|Esophagus|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C150-C155,C158-C159|Esophagus|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C150-C155,C158-C159|Esophagus|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C150-C155,C158-C159|Esophagus|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C150-C155,C158-C159|Esophagus|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C150-C155,C158-C159|Esophagus|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C150-C155,C158-C159|Esophagus|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C150-C155,C158-C159|Esophagus|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C150-C155,C158-C159|Esophagus|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C150-C155,C158-C159|Esophagus|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C150-C155,C158-C159|Esophagus|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C150-C155,C158-C159|Esophagus|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C150-C155,C158-C159|Esophagus|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C150-C155,C158-C159|Esophagus|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C150-C155,C158-C159|Esophagus|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8720/3|Melanoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8721/3|Nodular_Melanoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C150-C155,C158-C159|Esophagus|872|Melanoma|8723/3|Regressing_Melanoma
C150-C155,C158-C159|Esophagus|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C150-C155,C158-C159|Esophagus|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C150-C155,C158-C159|Esophagus|874|Nevus|8745/3|Desmoplastic_Melanoma
C150-C155,C158-C159|Esophagus|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C150-C155,C158-C159|Esophagus|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C150-C155,C158-C159|Esophagus|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C150-C155,C158-C159|Esophagus|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C150-C155,C158-C159|Esophagus|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C150-C155,C158-C159|Esophagus|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C150-C155,C158-C159|Esophagus|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C150-C155,C158-C159|Esophagus|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C150-C155,C158-C159|Esophagus|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C150-C155,C158-C159|Esophagus|898|Carcinosarcoma|8980/3|Carcinosarcoma
C150-C155,C158-C159|Esophagus|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C150-C155,C158-C159|Esophagus|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C150-C155,C158-C159|Esophagus|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C150-C155,C158-C159|Esophagus|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C150-C155,C158-C159|Esophagus|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C150-C155,C158-C159|Esophagus|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C150-C155,C158-C159|Esophagus|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C150-C155,C158-C159|Esophagus|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C150-C155,C158-C159|Esophagus|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C150-C155,C158-C159|Esophagus|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C150-C155,C158-C159|Esophagus|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C150-C155,C158-C159|Esophagus|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C150-C155,C158-C159|Esophagus|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C150-C155,C158-C159|Esophagus|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C150-C155,C158-C159|Esophagus|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C150-C155,C158-C159|Esophagus|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9731/3|Plasmacytoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C150-C155,C158-C159|Esophagus|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C150-C155,C158-C159|Esophagus|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C150-C155,C158-C159|Esophagus|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C150-C155,C158-C159|Esophagus|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C150-C155,C158-C159|Esophagus|975|Neoplasm|9750/3|Malignant_Histiocytosis
C150-C155,C158-C159|Esophagus|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C150-C155,C158-C159|Esophagus|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C150-C155,C158-C159|Esophagus|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C150-C155,C158-C159|Esophagus|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C150-C155,C158-C159|Esophagus|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C150-C155,C158-C159|Esophagus|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C150-C155,C158-C159|Esophagus|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C150-C155,C158-C159|Esophagus|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C150-C155,C158-C159|Esophagus|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C150-C155,C158-C159|Esophagus|981|Neoplasm|9812/3|Lymphoma
C150-C155,C158-C159|Esophagus|981|Neoplasm|9813/3|Lymphoma
C150-C155,C158-C159|Esophagus|981|Neoplasm|9814/3|Lymphoma
C150-C155,C158-C159|Esophagus|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C150-C155,C158-C159|Esophagus|981|Neoplasm|9816/3|Hypodiploid_ALL
C150-C155,C158-C159|Esophagus|981|Neoplasm|9817/3|Lymphoma
C150-C155,C158-C159|Esophagus|981|Neoplasm|9818/3|Lymphoma
C150-C155,C158-C159|Esophagus|981|Neoplasm|9819/3|Leukemia__B_Cell
C150-C155,C158-C159|Esophagus|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C150-C155,C158-C159|Esophagus|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C150-C155,C158-C159|Esophagus|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C150-C155,C158-C159|Esophagus|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C150-C155,C158-C159|Esophagus|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C150-C155,C158-C159|Esophagus|997|Neoplasm|9971/3|Polymorphic_PTLD
C150-C155,C158-C159|Esophagus|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C160-C166,C168-C169|Stomach|800|Neoplasm|8000/3|Malignant_Neoplasm
C160-C166,C168-C169|Stomach|800|Neoplasm|8001/3|Malignant_Cell
C160-C166,C168-C169|Stomach|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C160-C166,C168-C169|Stomach|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C160-C166,C168-C169|Stomach|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C160-C166,C168-C169|Stomach|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C160-C166,C168-C169|Stomach|801|Carcinoma|8010/2|In_Situ_Cancer
C160-C166,C168-C169|Stomach|801|Carcinoma|8010/3|Carcinoma
C160-C166,C168-C169|Stomach|801|Carcinoma|8011/3|Malignant_Epithelioma
C160-C166,C168-C169|Stomach|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C160-C166,C168-C169|Stomach|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C160-C166,C168-C169|Stomach|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C160-C166,C168-C169|Stomach|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C160-C166,C168-C169|Stomach|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C160-C166,C168-C169|Stomach|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C160-C166,C168-C169|Stomach|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C160-C166,C168-C169|Stomach|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C160-C166,C168-C169|Stomach|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C160-C166,C168-C169|Stomach|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C160-C166,C168-C169|Stomach|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C160-C166,C168-C169|Stomach|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C160-C166,C168-C169|Stomach|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C160-C166,C168-C169|Stomach|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C160-C166,C168-C169|Stomach|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C160-C166,C168-C169|Stomach|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C160-C166,C168-C169|Stomach|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C160-C166,C168-C169|Stomach|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C160-C166,C168-C169|Stomach|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C160-C166,C168-C169|Stomach|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C160-C166,C168-C169|Stomach|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8140/3|Adenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8142/3|Linitis_Plastica
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8144/3|Intestinal_Type_Adenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8145/3|Diffuse_Type_Adenocarcinoma
C160-C166,C168-C169|Stomach|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C160-C166,C168-C169|Stomach|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C160-C166,C168-C169|Stomach|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C160-C166,C168-C169|Stomach|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C160-C166,C168-C169|Stomach|821|Adenocarcinoma_In_Adenomatous_Polyp|8214/3|Gastric_Parietal_Cell_Adenocarcinoma
C160-C166,C168-C169|Stomach|822|Familial_Adenomatous_Polyposis|8220/2|Adenocarcinoma_In_Situ
C160-C166,C168-C169|Stomach|822|Familial_Adenomatous_Polyposis|8220/3|Familial_Adenomatous_Polyposis
C160-C166,C168-C169|Stomach|822|Familial_Adenomatous_Polyposis|8221/2|Adenomatous_Polyp
C160-C166,C168-C169|Stomach|822|Familial_Adenomatous_Polyposis|8221/3|Adenomatous_Polyp
C160-C166,C168-C169|Stomach|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C160-C166,C168-C169|Stomach|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C160-C166,C168-C169|Stomach|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C160-C166,C168-C169|Stomach|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C160-C166,C168-C169|Stomach|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C160-C166,C168-C169|Stomach|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C160-C166,C168-C169|Stomach|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C160-C166,C168-C169|Stomach|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C160-C166,C168-C169|Stomach|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C160-C166,C168-C169|Stomach|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C160-C166,C168-C169|Stomach|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C160-C166,C168-C169|Stomach|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C160-C166,C168-C169|Stomach|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C160-C166,C168-C169|Stomach|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C160-C166,C168-C169|Stomach|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C160-C166,C168-C169|Stomach|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C160-C166,C168-C169|Stomach|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C160-C166,C168-C169|Stomach|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C160-C166,C168-C169|Stomach|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C160-C166,C168-C169|Stomach|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C160-C166,C168-C169|Stomach|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C160-C166,C168-C169|Stomach|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C160-C166,C168-C169|Stomach|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C160-C166,C168-C169|Stomach|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C160-C166,C168-C169|Stomach|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C160-C166,C168-C169|Stomach|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C160-C166,C168-C169|Stomach|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C160-C166,C168-C169|Stomach|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C160-C166,C168-C169|Stomach|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C160-C166,C168-C169|Stomach|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C160-C166,C168-C169|Stomach|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C160-C166,C168-C169|Stomach|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8800/3|Sarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C160-C166,C168-C169|Stomach|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C160-C166,C168-C169|Stomach|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C160-C166,C168-C169|Stomach|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C160-C166,C168-C169|Stomach|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C160-C166,C168-C169|Stomach|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C160-C166,C168-C169|Stomach|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C160-C166,C168-C169|Stomach|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C160-C166,C168-C169|Stomach|893|Stromal_Sarcoma|8934/3|Carcinofibroma
C160-C166,C168-C169|Stomach|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C160-C166,C168-C169|Stomach|893|Stromal_Sarcoma|8936/3|High_Risk_Gastrointestinal_Stromal_Tumor
C160-C166,C168-C169|Stomach|898|Carcinosarcoma|8980/3|Carcinosarcoma
C160-C166,C168-C169|Stomach|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C160-C166,C168-C169|Stomach|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C160-C166,C168-C169|Stomach|959|Lymphoma|9590/3|Lymphoma
C160-C166,C168-C169|Stomach|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C160-C166,C168-C169|Stomach|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C160-C166,C168-C169|Stomach|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C160-C166,C168-C169|Stomach|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C160-C166,C168-C169|Stomach|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C160-C166,C168-C169|Stomach|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C160-C166,C168-C169|Stomach|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C160-C166,C168-C169|Stomach|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C160-C166,C168-C169|Stomach|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C160-C166,C168-C169|Stomach|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C160-C166,C168-C169|Stomach|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C160-C166,C168-C169|Stomach|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C160-C166,C168-C169|Stomach|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C160-C166,C168-C169|Stomach|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C160-C166,C168-C169|Stomach|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C160-C166,C168-C169|Stomach|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C160-C166,C168-C169|Stomach|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C160-C166,C168-C169|Stomach|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C160-C166,C168-C169|Stomach|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C160-C166,C168-C169|Stomach|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C160-C166,C168-C169|Stomach|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C160-C166,C168-C169|Stomach|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C160-C166,C168-C169|Stomach|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C160-C166,C168-C169|Stomach|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C160-C166,C168-C169|Stomach|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C160-C166,C168-C169|Stomach|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C160-C166,C168-C169|Stomach|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C160-C166,C168-C169|Stomach|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C160-C166,C168-C169|Stomach|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9731/3|Plasmacytoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9732/3|Plasma_Cell_Myeloma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C160-C166,C168-C169|Stomach|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C160-C166,C168-C169|Stomach|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C160-C166,C168-C169|Stomach|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C160-C166,C168-C169|Stomach|975|Neoplasm|9750/3|Malignant_Histiocytosis
C160-C166,C168-C169|Stomach|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C160-C166,C168-C169|Stomach|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C160-C166,C168-C169|Stomach|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C160-C166,C168-C169|Stomach|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C160-C166,C168-C169|Stomach|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C160-C166,C168-C169|Stomach|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C160-C166,C168-C169|Stomach|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C160-C166,C168-C169|Stomach|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C160-C166,C168-C169|Stomach|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C160-C166,C168-C169|Stomach|981|Neoplasm|9812/3|Lymphoma
C160-C166,C168-C169|Stomach|981|Neoplasm|9813/3|Lymphoma
C160-C166,C168-C169|Stomach|981|Neoplasm|9814/3|Lymphoma
C160-C166,C168-C169|Stomach|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C160-C166,C168-C169|Stomach|981|Neoplasm|9816/3|Hypodiploid_ALL
C160-C166,C168-C169|Stomach|981|Neoplasm|9817/3|Lymphoma
C160-C166,C168-C169|Stomach|981|Neoplasm|9818/3|Lymphoma
C160-C166,C168-C169|Stomach|981|Neoplasm|9819/3|Leukemia__B_Cell
C160-C166,C168-C169|Stomach|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C160-C166,C168-C169|Stomach|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C160-C166,C168-C169|Stomach|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C160-C166,C168-C169|Stomach|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C160-C166,C168-C169|Stomach|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C160-C166,C168-C169|Stomach|997|Neoplasm|9971/3|Polymorphic_PTLD
C160-C166,C168-C169|Stomach|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C170-C173,C178-C179|Small_Intestine|800|Neoplasm|8000/3|Malignant_Neoplasm
C170-C173,C178-C179|Small_Intestine|800|Neoplasm|8001/3|Malignant_Cell
C170-C173,C178-C179|Small_Intestine|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C170-C173,C178-C179|Small_Intestine|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C170-C173,C178-C179|Small_Intestine|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C170-C173,C178-C179|Small_Intestine|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C170-C173,C178-C179|Small_Intestine|801|Carcinoma|8010/2|In_Situ_Cancer
C170-C173,C178-C179|Small_Intestine|801|Carcinoma|8010/3|Carcinoma
C170-C173,C178-C179|Small_Intestine|801|Carcinoma|8011/3|Malignant_Epithelioma
C170-C173,C178-C179|Small_Intestine|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C170-C173,C178-C179|Small_Intestine|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C170-C173,C178-C179|Small_Intestine|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C170-C173,C178-C179|Small_Intestine|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C170-C173,C178-C179|Small_Intestine|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C170-C173,C178-C179|Small_Intestine|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C170-C173,C178-C179|Small_Intestine|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C170-C173,C178-C179|Small_Intestine|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C170-C173,C178-C179|Small_Intestine|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C170-C173,C178-C179|Small_Intestine|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C170-C173,C178-C179|Small_Intestine|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C170-C173,C178-C179|Small_Intestine|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C170-C173,C178-C179|Small_Intestine|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C170-C173,C178-C179|Small_Intestine|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C170-C173,C178-C179|Small_Intestine|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C170-C173,C178-C179|Small_Intestine|814|Adenocarcinoma|8140/3|Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|814|Adenocarcinoma|8145/3|Diffuse_Type_Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C170-C173,C178-C179|Small_Intestine|815|Endocrine_Gland_Neoplasms|8152/3|Malignant_Pancreatic_Glucagonoma
C170-C173,C178-C179|Small_Intestine|815|Endocrine_Gland_Neoplasms|8153/3|Malignant_Gastrinoma
C170-C173,C178-C179|Small_Intestine|815|Endocrine_Gland_Neoplasms|8156/3|Malignant_Somatostatinoma
C170-C173,C178-C179|Small_Intestine|815|Endocrine_Gland_Neoplasms|8157/3|Malignant_Enteroglucagonoma
C170-C173,C178-C179|Small_Intestine|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C170-C173,C178-C179|Small_Intestine|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C170-C173,C178-C179|Small_Intestine|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C170-C173,C178-C179|Small_Intestine|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C170-C173,C178-C179|Small_Intestine|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C170-C173,C178-C179|Small_Intestine|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C170-C173,C178-C179|Small_Intestine|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C170-C173,C178-C179|Small_Intestine|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C170-C173,C178-C179|Small_Intestine|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C170-C173,C178-C179|Small_Intestine|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C170-C173,C178-C179|Small_Intestine|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C170-C173,C178-C179|Small_Intestine|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C170-C173,C178-C179|Small_Intestine|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C170-C173,C178-C179|Small_Intestine|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C170-C173,C178-C179|Small_Intestine|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C170-C173,C178-C179|Small_Intestine|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C170-C173,C178-C179|Small_Intestine|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C170-C173,C178-C179|Small_Intestine|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C170-C173,C178-C179|Small_Intestine|871|Malignant_Glomus_Tumor|8710/3|Malignant_Glomus_Tumor
C170-C173,C178-C179|Small_Intestine|880|Sarcoma|8800/3|Sarcoma
C170-C173,C178-C179|Small_Intestine|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C170-C173,C178-C179|Small_Intestine|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C170-C173,C178-C179|Small_Intestine|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C170-C173,C178-C179|Small_Intestine|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C170-C173,C178-C179|Small_Intestine|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C170-C173,C178-C179|Small_Intestine|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C170-C173,C178-C179|Small_Intestine|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C170-C173,C178-C179|Small_Intestine|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C170-C173,C178-C179|Small_Intestine|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C170-C173,C178-C179|Small_Intestine|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C170-C173,C178-C179|Small_Intestine|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C170-C173,C178-C179|Small_Intestine|882|Sarcoma|8825/3|Sarcoma
C170-C173,C178-C179|Small_Intestine|885|Liposarcoma|8850/3|Liposarcoma
C170-C173,C178-C179|Small_Intestine|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C170-C173,C178-C179|Small_Intestine|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C170-C173,C178-C179|Small_Intestine|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C170-C173,C178-C179|Small_Intestine|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C170-C173,C178-C179|Small_Intestine|885|Liposarcoma|8855/3|Liposarcoma
C170-C173,C178-C179|Small_Intestine|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C170-C173,C178-C179|Small_Intestine|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C170-C173,C178-C179|Small_Intestine|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C170-C173,C178-C179|Small_Intestine|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C170-C173,C178-C179|Small_Intestine|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C170-C173,C178-C179|Small_Intestine|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C170-C173,C178-C179|Small_Intestine|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C170-C173,C178-C179|Small_Intestine|893|Stromal_Sarcoma|8934/3|Carcinofibroma
C170-C173,C178-C179|Small_Intestine|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C170-C173,C178-C179|Small_Intestine|893|Stromal_Sarcoma|8936/3|High_Risk_Gastrointestinal_Stromal_Tumor
C170-C173,C178-C179|Small_Intestine|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C170-C173,C178-C179|Small_Intestine|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C170-C173,C178-C179|Small_Intestine|959|Lymphoma|9590/3|Lymphoma
C170-C173,C178-C179|Small_Intestine|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C170-C173,C178-C179|Small_Intestine|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C170-C173,C178-C179|Small_Intestine|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C170-C173,C178-C179|Small_Intestine|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C170-C173,C178-C179|Small_Intestine|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C170-C173,C178-C179|Small_Intestine|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C170-C173,C178-C179|Small_Intestine|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C170-C173,C178-C179|Small_Intestine|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C170-C173,C178-C179|Small_Intestine|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C170-C173,C178-C179|Small_Intestine|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C170-C173,C178-C179|Small_Intestine|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C170-C173,C178-C179|Small_Intestine|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C170-C173,C178-C179|Small_Intestine|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C170-C173,C178-C179|Small_Intestine|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C170-C173,C178-C179|Small_Intestine|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C170-C173,C178-C179|Small_Intestine|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C170-C173,C178-C179|Small_Intestine|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C170-C173,C178-C179|Small_Intestine|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C170-C173,C178-C179|Small_Intestine|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C170-C173,C178-C179|Small_Intestine|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C170-C173,C178-C179|Small_Intestine|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C170-C173,C178-C179|Small_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C170-C173,C178-C179|Small_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C170-C173,C178-C179|Small_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C170-C173,C178-C179|Small_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C170-C173,C178-C179|Small_Intestine|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C170-C173,C178-C179|Small_Intestine|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C170-C173,C178-C179|Small_Intestine|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C170-C173,C178-C179|Small_Intestine|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C170-C173,C178-C179|Small_Intestine|973|Plasmacytoma|9731/3|Plasmacytoma
C170-C173,C178-C179|Small_Intestine|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C170-C173,C178-C179|Small_Intestine|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C170-C173,C178-C179|Small_Intestine|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C170-C173,C178-C179|Small_Intestine|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C170-C173,C178-C179|Small_Intestine|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C170-C173,C178-C179|Small_Intestine|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C170-C173,C178-C179|Small_Intestine|975|Neoplasm|9750/3|Malignant_Histiocytosis
C170-C173,C178-C179|Small_Intestine|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C170-C173,C178-C179|Small_Intestine|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C170-C173,C178-C179|Small_Intestine|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C170-C173,C178-C179|Small_Intestine|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C170-C173,C178-C179|Small_Intestine|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C170-C173,C178-C179|Small_Intestine|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C170-C173,C178-C179|Small_Intestine|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C170-C173,C178-C179|Small_Intestine|976|Immunoproliferative_Disorder|9764/3|Immunoproliferative_Disorder
C170-C173,C178-C179|Small_Intestine|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9812/3|Lymphoma
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9813/3|Lymphoma
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9814/3|Lymphoma
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9816/3|Hypodiploid_ALL
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9817/3|Lymphoma
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9818/3|Lymphoma
C170-C173,C178-C179|Small_Intestine|981|Neoplasm|9819/3|Leukemia__B_Cell
C170-C173,C178-C179|Small_Intestine|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C170-C173,C178-C179|Small_Intestine|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C170-C173,C178-C179|Small_Intestine|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C170-C173,C178-C179|Small_Intestine|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C170-C173,C178-C179|Small_Intestine|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C170-C173,C178-C179|Small_Intestine|997|Neoplasm|9971/3|Polymorphic_PTLD
C170-C173,C178-C179|Small_Intestine|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C180, C182-C189, C199|Large_Intestine|800|Neoplasm|8000/3|Malignant_Neoplasm
C180, C182-C189, C199|Large_Intestine|800|Neoplasm|8001/3|Malignant_Cell
C180, C182-C189, C199|Large_Intestine|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C180, C182-C189, C199|Large_Intestine|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C180, C182-C189, C199|Large_Intestine|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C180, C182-C189, C199|Large_Intestine|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C180, C182-C189, C199|Large_Intestine|801|Carcinoma|8010/2|In_Situ_Cancer
C180, C182-C189, C199|Large_Intestine|801|Carcinoma|8010/3|Carcinoma
C180, C182-C189, C199|Large_Intestine|801|Carcinoma|8011/3|Malignant_Epithelioma
C180, C182-C189, C199|Large_Intestine|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C180, C182-C189, C199|Large_Intestine|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C180, C182-C189, C199|Large_Intestine|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C180, C182-C189, C199|Large_Intestine|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C180, C182-C189, C199|Large_Intestine|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C180, C182-C189, C199|Large_Intestine|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C180, C182-C189, C199|Large_Intestine|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C180, C182-C189, C199|Large_Intestine|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C180, C182-C189, C199|Large_Intestine|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C180, C182-C189, C199|Large_Intestine|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C180, C182-C189, C199|Large_Intestine|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C180, C182-C189, C199|Large_Intestine|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C180, C182-C189, C199|Large_Intestine|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C180, C182-C189, C199|Large_Intestine|814|Adenocarcinoma|8140/3|Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|814|Adenocarcinoma|8145/3|Diffuse_Type_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C180, C182-C189, C199|Large_Intestine|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C180, C182-C189, C199|Large_Intestine|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C180, C182-C189, C199|Large_Intestine|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|821|Adenocarcinoma_In_Adenomatous_Polyp|8213/3|Serrated_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|822|Familial_Adenomatous_Polyposis|8220/2|Adenocarcinoma_In_Situ
C180, C182-C189, C199|Large_Intestine|822|Familial_Adenomatous_Polyposis|8220/3|Familial_Adenomatous_Polyposis
C180, C182-C189, C199|Large_Intestine|822|Familial_Adenomatous_Polyposis|8221/2|Adenomatous_Polyp
C180, C182-C189, C199|Large_Intestine|822|Familial_Adenomatous_Polyposis|8221/3|Adenomatous_Polyp
C180, C182-C189, C199|Large_Intestine|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C180, C182-C189, C199|Large_Intestine|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C180, C182-C189, C199|Large_Intestine|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C180, C182-C189, C199|Large_Intestine|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C180, C182-C189, C199|Large_Intestine|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C180, C182-C189, C199|Large_Intestine|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C180, C182-C189, C199|Large_Intestine|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C180, C182-C189, C199|Large_Intestine|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C180, C182-C189, C199|Large_Intestine|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C180, C182-C189, C199|Large_Intestine|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C180, C182-C189, C199|Large_Intestine|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C180, C182-C189, C199|Large_Intestine|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C180, C182-C189, C199|Large_Intestine|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C180, C182-C189, C199|Large_Intestine|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C180, C182-C189, C199|Large_Intestine|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C180, C182-C189, C199|Large_Intestine|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C180, C182-C189, C199|Large_Intestine|826|Papillary_Adenocarcinoma|8265/3|Micropapillary_Carcinoma
C180, C182-C189, C199|Large_Intestine|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C180, C182-C189, C199|Large_Intestine|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C180, C182-C189, C199|Large_Intestine|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C180, C182-C189, C199|Large_Intestine|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C180, C182-C189, C199|Large_Intestine|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C180, C182-C189, C199|Large_Intestine|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C180, C182-C189, C199|Large_Intestine|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C180, C182-C189, C199|Large_Intestine|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C180, C182-C189, C199|Large_Intestine|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C180, C182-C189, C199|Large_Intestine|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C180, C182-C189, C199|Large_Intestine|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C180, C182-C189, C199|Large_Intestine|880|Sarcoma|8800/3|Sarcoma
C180, C182-C189, C199|Large_Intestine|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C180, C182-C189, C199|Large_Intestine|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C180, C182-C189, C199|Large_Intestine|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C180, C182-C189, C199|Large_Intestine|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C180, C182-C189, C199|Large_Intestine|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C180, C182-C189, C199|Large_Intestine|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C180, C182-C189, C199|Large_Intestine|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C180, C182-C189, C199|Large_Intestine|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C180, C182-C189, C199|Large_Intestine|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C180, C182-C189, C199|Large_Intestine|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C180, C182-C189, C199|Large_Intestine|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C180, C182-C189, C199|Large_Intestine|882|Sarcoma|8825/3|Sarcoma
C180, C182-C189, C199|Large_Intestine|885|Liposarcoma|8850/3|Liposarcoma
C180, C182-C189, C199|Large_Intestine|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C180, C182-C189, C199|Large_Intestine|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C180, C182-C189, C199|Large_Intestine|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C180, C182-C189, C199|Large_Intestine|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C180, C182-C189, C199|Large_Intestine|885|Liposarcoma|8855/3|Liposarcoma
C180, C182-C189, C199|Large_Intestine|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C180, C182-C189, C199|Large_Intestine|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C180, C182-C189, C199|Large_Intestine|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C180, C182-C189, C199|Large_Intestine|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C180, C182-C189, C199|Large_Intestine|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C180, C182-C189, C199|Large_Intestine|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C180, C182-C189, C199|Large_Intestine|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C180, C182-C189, C199|Large_Intestine|893|Stromal_Sarcoma|8934/3|Carcinofibroma
C180, C182-C189, C199|Large_Intestine|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C180, C182-C189, C199|Large_Intestine|893|Stromal_Sarcoma|8936/3|High_Risk_Gastrointestinal_Stromal_Tumor
C180, C182-C189, C199|Large_Intestine|898|Carcinosarcoma|8980/3|Carcinosarcoma
C180, C182-C189, C199|Large_Intestine|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C180, C182-C189, C199|Large_Intestine|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C180, C182-C189, C199|Large_Intestine|959|Lymphoma|9590/3|Lymphoma
C180, C182-C189, C199|Large_Intestine|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C180, C182-C189, C199|Large_Intestine|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C180, C182-C189, C199|Large_Intestine|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C180, C182-C189, C199|Large_Intestine|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C180, C182-C189, C199|Large_Intestine|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C180, C182-C189, C199|Large_Intestine|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C180, C182-C189, C199|Large_Intestine|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C180, C182-C189, C199|Large_Intestine|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C180, C182-C189, C199|Large_Intestine|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C180, C182-C189, C199|Large_Intestine|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C180, C182-C189, C199|Large_Intestine|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C180, C182-C189, C199|Large_Intestine|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C180, C182-C189, C199|Large_Intestine|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C180, C182-C189, C199|Large_Intestine|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C180, C182-C189, C199|Large_Intestine|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C180, C182-C189, C199|Large_Intestine|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C180, C182-C189, C199|Large_Intestine|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C180, C182-C189, C199|Large_Intestine|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C180, C182-C189, C199|Large_Intestine|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C180, C182-C189, C199|Large_Intestine|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C180, C182-C189, C199|Large_Intestine|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C180, C182-C189, C199|Large_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C180, C182-C189, C199|Large_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C180, C182-C189, C199|Large_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C180, C182-C189, C199|Large_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C180, C182-C189, C199|Large_Intestine|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C180, C182-C189, C199|Large_Intestine|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C180, C182-C189, C199|Large_Intestine|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C180, C182-C189, C199|Large_Intestine|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C180, C182-C189, C199|Large_Intestine|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C180, C182-C189, C199|Large_Intestine|973|Plasmacytoma|9731/3|Plasmacytoma
C180, C182-C189, C199|Large_Intestine|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C180, C182-C189, C199|Large_Intestine|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C180, C182-C189, C199|Large_Intestine|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C180, C182-C189, C199|Large_Intestine|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C180, C182-C189, C199|Large_Intestine|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C180, C182-C189, C199|Large_Intestine|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C180, C182-C189, C199|Large_Intestine|975|Neoplasm|9750/3|Malignant_Histiocytosis
C180, C182-C189, C199|Large_Intestine|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C180, C182-C189, C199|Large_Intestine|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C180, C182-C189, C199|Large_Intestine|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C180, C182-C189, C199|Large_Intestine|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C180, C182-C189, C199|Large_Intestine|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C180, C182-C189, C199|Large_Intestine|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C180, C182-C189, C199|Large_Intestine|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C180, C182-C189, C199|Large_Intestine|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9812/3|Lymphoma
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9813/3|Lymphoma
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9814/3|Lymphoma
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9816/3|Hypodiploid_ALL
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9817/3|Lymphoma
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9818/3|Lymphoma
C180, C182-C189, C199|Large_Intestine|981|Neoplasm|9819/3|Leukemia__B_Cell
C180, C182-C189, C199|Large_Intestine|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C180, C182-C189, C199|Large_Intestine|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C180, C182-C189, C199|Large_Intestine|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C180, C182-C189, C199|Large_Intestine|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C180, C182-C189, C199|Large_Intestine|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C180, C182-C189, C199|Large_Intestine|997|Neoplasm|9971/3|Polymorphic_PTLD
C180, C182-C189, C199|Large_Intestine|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C181|Appendix|800|Neoplasm|8000/3|Malignant_Neoplasm
C181|Appendix|800|Neoplasm|8001/3|Malignant_Cell
C181|Appendix|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C181|Appendix|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C181|Appendix|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C181|Appendix|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C181|Appendix|801|Carcinoma|8010/2|In_Situ_Cancer
C181|Appendix|801|Carcinoma|8010/3|Carcinoma
C181|Appendix|801|Carcinoma|8011/3|Malignant_Epithelioma
C181|Appendix|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C181|Appendix|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C181|Appendix|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C181|Appendix|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C181|Appendix|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C181|Appendix|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C181|Appendix|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C181|Appendix|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C181|Appendix|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C181|Appendix|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C181|Appendix|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C181|Appendix|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C181|Appendix|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C181|Appendix|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C181|Appendix|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C181|Appendix|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C181|Appendix|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C181|Appendix|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C181|Appendix|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C181|Appendix|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C181|Appendix|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C181|Appendix|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C181|Appendix|814|Adenocarcinoma|8140/3|Adenocarcinoma
C181|Appendix|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C181|Appendix|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C181|Appendix|814|Adenocarcinoma|8145/3|Diffuse_Type_Adenocarcinoma
C181|Appendix|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C181|Appendix|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C181|Appendix|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C181|Appendix|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C181|Appendix|822|Familial_Adenomatous_Polyposis|8220/2|Adenocarcinoma_In_Situ
C181|Appendix|822|Familial_Adenomatous_Polyposis|8220/3|Familial_Adenomatous_Polyposis
C181|Appendix|822|Familial_Adenomatous_Polyposis|8221/2|Adenomatous_Polyp
C181|Appendix|822|Familial_Adenomatous_Polyposis|8221/3|Adenomatous_Polyp
C181|Appendix|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C181|Appendix|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C181|Appendix|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C181|Appendix|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C181|Appendix|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C181|Appendix|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C181|Appendix|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C181|Appendix|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C181|Appendix|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C181|Appendix|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C181|Appendix|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C181|Appendix|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C181|Appendix|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C181|Appendix|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C181|Appendix|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C181|Appendix|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C181|Appendix|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C181|Appendix|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C181|Appendix|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C181|Appendix|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C181|Appendix|847|Mucinous_Cystadenocarcinoma|8470/2|Mucinous_Cystadenocarcinoma
C181|Appendix|847|Mucinous_Cystadenocarcinoma|8470/3|Mucinous_Cystadenocarcinoma
C181|Appendix|847|Mucinous_Cystadenocarcinoma|8471/3|Papillary_Mucinous_Cystadenocarcinoma
C181|Appendix|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C181|Appendix|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C181|Appendix|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C181|Appendix|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C181|Appendix|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C181|Appendix|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C181|Appendix|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C181|Appendix|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C181|Appendix|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C181|Appendix|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C181|Appendix|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C181|Appendix|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C181|Appendix|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C181|Appendix|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C181|Appendix|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C181|Appendix|880|Sarcoma|8800/3|Sarcoma
C181|Appendix|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C181|Appendix|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C181|Appendix|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C181|Appendix|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C181|Appendix|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C181|Appendix|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C181|Appendix|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C181|Appendix|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C181|Appendix|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C181|Appendix|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C181|Appendix|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C181|Appendix|882|Sarcoma|8825/3|Sarcoma
C181|Appendix|885|Liposarcoma|8850/3|Liposarcoma
C181|Appendix|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C181|Appendix|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C181|Appendix|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C181|Appendix|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C181|Appendix|885|Liposarcoma|8855/3|Liposarcoma
C181|Appendix|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C181|Appendix|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C181|Appendix|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C181|Appendix|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C181|Appendix|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C181|Appendix|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C181|Appendix|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C181|Appendix|893|Stromal_Sarcoma|8934/3|Carcinofibroma
C181|Appendix|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C181|Appendix|893|Stromal_Sarcoma|8936/3|High_Risk_Gastrointestinal_Stromal_Tumor
C181|Appendix|898|Carcinosarcoma|8980/3|Carcinosarcoma
C181|Appendix|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C181|Appendix|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C181|Appendix|959|Lymphoma|9590/3|Lymphoma
C181|Appendix|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C181|Appendix|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C181|Appendix|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C181|Appendix|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C181|Appendix|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C181|Appendix|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C181|Appendix|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C181|Appendix|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C181|Appendix|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C181|Appendix|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C181|Appendix|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C181|Appendix|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C181|Appendix|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C181|Appendix|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C181|Appendix|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C181|Appendix|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C181|Appendix|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C181|Appendix|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C181|Appendix|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C181|Appendix|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C181|Appendix|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C181|Appendix|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C181|Appendix|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C181|Appendix|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C181|Appendix|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C181|Appendix|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C181|Appendix|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C181|Appendix|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C181|Appendix|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C181|Appendix|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C181|Appendix|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C181|Appendix|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C181|Appendix|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C181|Appendix|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C181|Appendix|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C181|Appendix|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C181|Appendix|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C181|Appendix|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C181|Appendix|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C181|Appendix|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C181|Appendix|973|Plasmacytoma|9731/3|Plasmacytoma
C181|Appendix|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C181|Appendix|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C181|Appendix|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C181|Appendix|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C181|Appendix|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C181|Appendix|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C181|Appendix|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C181|Appendix|975|Neoplasm|9750/3|Malignant_Histiocytosis
C181|Appendix|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C181|Appendix|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C181|Appendix|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C181|Appendix|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C181|Appendix|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C181|Appendix|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C181|Appendix|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C181|Appendix|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C181|Appendix|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C181|Appendix|981|Neoplasm|9812/3|Lymphoma
C181|Appendix|981|Neoplasm|9813/3|Lymphoma
C181|Appendix|981|Neoplasm|9814/3|Lymphoma
C181|Appendix|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C181|Appendix|981|Neoplasm|9816/3|Hypodiploid_ALL
C181|Appendix|981|Neoplasm|9817/3|Lymphoma
C181|Appendix|981|Neoplasm|9818/3|Lymphoma
C181|Appendix|981|Neoplasm|9819/3|Leukemia__B_Cell
C181|Appendix|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C181|Appendix|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C181|Appendix|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C181|Appendix|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C181|Appendix|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C181|Appendix|997|Neoplasm|9971/3|Polymorphic_PTLD
C181|Appendix|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C209|Rectal|800|Neoplasm|8000/3|Malignant_Neoplasm
C209|Rectal|800|Neoplasm|8001/3|Malignant_Cell
C209|Rectal|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C209|Rectal|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C209|Rectal|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C209|Rectal|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C209|Rectal|801|Carcinoma|8010/2|In_Situ_Cancer
C209|Rectal|801|Carcinoma|8010/3|Carcinoma
C209|Rectal|801|Carcinoma|8011/3|Malignant_Epithelioma
C209|Rectal|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C209|Rectal|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C209|Rectal|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C209|Rectal|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C209|Rectal|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C209|Rectal|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C209|Rectal|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C209|Rectal|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C209|Rectal|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C209|Rectal|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C209|Rectal|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C209|Rectal|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C209|Rectal|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C209|Rectal|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C209|Rectal|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C209|Rectal|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C209|Rectal|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C209|Rectal|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C209|Rectal|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C209|Rectal|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C209|Rectal|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C209|Rectal|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C209|Rectal|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C209|Rectal|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C209|Rectal|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C209|Rectal|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C209|Rectal|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C209|Rectal|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C209|Rectal|814|Adenocarcinoma|8140/3|Adenocarcinoma
C209|Rectal|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C209|Rectal|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C209|Rectal|814|Adenocarcinoma|8145/3|Diffuse_Type_Adenocarcinoma
C209|Rectal|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C209|Rectal|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C209|Rectal|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C209|Rectal|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C209|Rectal|821|Adenocarcinoma_In_Adenomatous_Polyp|8213/3|Serrated_Adenocarcinoma
C209|Rectal|822|Familial_Adenomatous_Polyposis|8220/2|Adenocarcinoma_In_Situ
C209|Rectal|822|Familial_Adenomatous_Polyposis|8220/3|Familial_Adenomatous_Polyposis
C209|Rectal|822|Familial_Adenomatous_Polyposis|8221/2|Adenomatous_Polyp
C209|Rectal|822|Familial_Adenomatous_Polyposis|8221/3|Adenomatous_Polyp
C209|Rectal|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C209|Rectal|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C209|Rectal|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C209|Rectal|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C209|Rectal|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C209|Rectal|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C209|Rectal|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C209|Rectal|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C209|Rectal|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C209|Rectal|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C209|Rectal|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C209|Rectal|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C209|Rectal|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C209|Rectal|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C209|Rectal|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C209|Rectal|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C209|Rectal|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C209|Rectal|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C209|Rectal|826|Papillary_Adenocarcinoma|8265/3|Micropapillary_Carcinoma
C209|Rectal|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C209|Rectal|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C209|Rectal|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C209|Rectal|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C209|Rectal|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C209|Rectal|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C209|Rectal|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C209|Rectal|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C209|Rectal|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C209|Rectal|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C209|Rectal|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C209|Rectal|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C209|Rectal|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C209|Rectal|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C209|Rectal|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C209|Rectal|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C209|Rectal|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C209|Rectal|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C209|Rectal|872|Melanoma|8720/3|Melanoma
C209|Rectal|872|Melanoma|8721/3|Nodular_Melanoma
C209|Rectal|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C209|Rectal|872|Melanoma|8723/3|Regressing_Melanoma
C209|Rectal|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C209|Rectal|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C209|Rectal|874|Nevus|8745/3|Desmoplastic_Melanoma
C209|Rectal|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C209|Rectal|876|Nevus|8761/3|Giant_Congenital_Nevus
C209|Rectal|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C209|Rectal|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C209|Rectal|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C209|Rectal|880|Sarcoma|8800/3|Sarcoma
C209|Rectal|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C209|Rectal|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C209|Rectal|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C209|Rectal|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C209|Rectal|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C209|Rectal|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C209|Rectal|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C209|Rectal|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C209|Rectal|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C209|Rectal|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C209|Rectal|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C209|Rectal|882|Sarcoma|8825/3|Sarcoma
C209|Rectal|885|Liposarcoma|8850/3|Liposarcoma
C209|Rectal|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C209|Rectal|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C209|Rectal|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C209|Rectal|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C209|Rectal|885|Liposarcoma|8855/3|Liposarcoma
C209|Rectal|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C209|Rectal|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C209|Rectal|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C209|Rectal|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C209|Rectal|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C209|Rectal|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C209|Rectal|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C209|Rectal|893|Stromal_Sarcoma|8934/3|Carcinofibroma
C209|Rectal|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C209|Rectal|893|Stromal_Sarcoma|8936/3|High_Risk_Gastrointestinal_Stromal_Tumor
C209|Rectal|898|Carcinosarcoma|8980/3|Carcinosarcoma
C209|Rectal|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C209|Rectal|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C209|Rectal|959|Lymphoma|9590/3|Lymphoma
C209|Rectal|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C209|Rectal|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C209|Rectal|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C209|Rectal|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C209|Rectal|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C209|Rectal|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C209|Rectal|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C209|Rectal|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C209|Rectal|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C209|Rectal|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C209|Rectal|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C209|Rectal|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C209|Rectal|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C209|Rectal|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C209|Rectal|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C209|Rectal|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C209|Rectal|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C209|Rectal|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C209|Rectal|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C209|Rectal|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C209|Rectal|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C209|Rectal|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C209|Rectal|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C209|Rectal|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C209|Rectal|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C209|Rectal|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C209|Rectal|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C209|Rectal|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C209|Rectal|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C209|Rectal|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C209|Rectal|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C209|Rectal|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C209|Rectal|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C209|Rectal|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C209|Rectal|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C209|Rectal|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C209|Rectal|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C209|Rectal|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C209|Rectal|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C209|Rectal|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C209|Rectal|973|Plasmacytoma|9731/3|Plasmacytoma
C209|Rectal|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C209|Rectal|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C209|Rectal|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C209|Rectal|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C209|Rectal|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C209|Rectal|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C209|Rectal|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C209|Rectal|975|Neoplasm|9750/3|Malignant_Histiocytosis
C209|Rectal|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C209|Rectal|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C209|Rectal|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C209|Rectal|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C209|Rectal|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C209|Rectal|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C209|Rectal|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C209|Rectal|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C209|Rectal|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C209|Rectal|981|Neoplasm|9812/3|Lymphoma
C209|Rectal|981|Neoplasm|9813/3|Lymphoma
C209|Rectal|981|Neoplasm|9814/3|Lymphoma
C209|Rectal|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C209|Rectal|981|Neoplasm|9816/3|Hypodiploid_ALL
C209|Rectal|981|Neoplasm|9817/3|Lymphoma
C209|Rectal|981|Neoplasm|9818/3|Lymphoma
C209|Rectal|981|Neoplasm|9819/3|Leukemia__B_Cell
C209|Rectal|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C209|Rectal|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C209|Rectal|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C209|Rectal|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C209|Rectal|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C209|Rectal|997|Neoplasm|9971/3|Polymorphic_PTLD
C209|Rectal|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C210-C212,C218|Anal_Canal|800|Neoplasm|8000/3|Malignant_Neoplasm
C210-C212,C218|Anal_Canal|800|Neoplasm|8001/3|Malignant_Cell
C210-C212,C218|Anal_Canal|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C210-C212,C218|Anal_Canal|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C210-C212,C218|Anal_Canal|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C210-C212,C218|Anal_Canal|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C210-C212,C218|Anal_Canal|801|Carcinoma|8010/2|In_Situ_Cancer
C210-C212,C218|Anal_Canal|801|Carcinoma|8010/3|Carcinoma
C210-C212,C218|Anal_Canal|801|Carcinoma|8011/3|Malignant_Epithelioma
C210-C212,C218|Anal_Canal|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C210-C212,C218|Anal_Canal|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C210-C212,C218|Anal_Canal|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C210-C212,C218|Anal_Canal|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C210-C212,C218|Anal_Canal|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C210-C212,C218|Anal_Canal|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C210-C212,C218|Anal_Canal|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C210-C212,C218|Anal_Canal|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C210-C212,C218|Anal_Canal|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C210-C212,C218|Anal_Canal|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C210-C212,C218|Anal_Canal|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C210-C212,C218|Anal_Canal|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C210-C212,C218|Anal_Canal|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C210-C212,C218|Anal_Canal|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8077/2|Intraepithelial_Neoplasia
C210-C212,C218|Anal_Canal|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C210-C212,C218|Anal_Canal|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C210-C212,C218|Anal_Canal|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C210-C212,C218|Anal_Canal|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C210-C212,C218|Anal_Canal|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C210-C212,C218|Anal_Canal|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C210-C212,C218|Anal_Canal|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C210-C212,C218|Anal_Canal|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C210-C212,C218|Anal_Canal|814|Adenocarcinoma|8140/3|Adenocarcinoma
C210-C212,C218|Anal_Canal|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C210-C212,C218|Anal_Canal|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C210-C212,C218|Anal_Canal|814|Adenocarcinoma|8145/3|Diffuse_Type_Adenocarcinoma
C210-C212,C218|Anal_Canal|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C210-C212,C218|Anal_Canal|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C210-C212,C218|Anal_Canal|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C210-C212,C218|Anal_Canal|821|Adenocarcinoma_In_Adenomatous_Polyp|8215/3|Anal_Glands_Adenocarcinoma
C210-C212,C218|Anal_Canal|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C210-C212,C218|Anal_Canal|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C210-C212,C218|Anal_Canal|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C210-C212,C218|Anal_Canal|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C210-C212,C218|Anal_Canal|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C210-C212,C218|Anal_Canal|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C210-C212,C218|Anal_Canal|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C210-C212,C218|Anal_Canal|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C210-C212,C218|Anal_Canal|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C210-C212,C218|Anal_Canal|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C210-C212,C218|Anal_Canal|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C210-C212,C218|Anal_Canal|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C210-C212,C218|Anal_Canal|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C210-C212,C218|Anal_Canal|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C210-C212,C218|Anal_Canal|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C210-C212,C218|Anal_Canal|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C210-C212,C218|Anal_Canal|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C210-C212,C218|Anal_Canal|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C210-C212,C218|Anal_Canal|850|Ductal_Carcinoma|8500/2|Ductal_Breast_Carcinoma_In_Situ
C210-C212,C218|Anal_Canal|850|Ductal_Carcinoma|8500/3|Invasive_Carcinoma
C210-C212,C218|Anal_Canal|850|Ductal_Carcinoma|8503/2|Intraductal_Papillary_Breast_Carcinoma
C210-C212,C218|Anal_Canal|850|Ductal_Carcinoma|8503/3|Intraductal_Papillary_Breast_Carcinoma
C210-C212,C218|Anal_Canal|850|Ductal_Carcinoma|8504/2|Intracystic_Papillary_Breast_Carcinoma
C210-C212,C218|Anal_Canal|850|Ductal_Carcinoma|8504/3|Intracystic_Papillary_Breast_Carcinoma
C210-C212,C218|Anal_Canal|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C210-C212,C218|Anal_Canal|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C210-C212,C218|Anal_Canal|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C210-C212,C218|Anal_Canal|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C210-C212,C218|Anal_Canal|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C210-C212,C218|Anal_Canal|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C210-C212,C218|Anal_Canal|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C210-C212,C218|Anal_Canal|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C210-C212,C218|Anal_Canal|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C210-C212,C218|Anal_Canal|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C210-C212,C218|Anal_Canal|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C210-C212,C218|Anal_Canal|872|Melanoma|8720/3|Melanoma
C210-C212,C218|Anal_Canal|872|Melanoma|8721/3|Nodular_Melanoma
C210-C212,C218|Anal_Canal|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C210-C212,C218|Anal_Canal|872|Melanoma|8723/3|Regressing_Melanoma
C210-C212,C218|Anal_Canal|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C210-C212,C218|Anal_Canal|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C210-C212,C218|Anal_Canal|874|Nevus|8745/3|Desmoplastic_Melanoma
C210-C212,C218|Anal_Canal|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C210-C212,C218|Anal_Canal|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C210-C212,C218|Anal_Canal|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C210-C212,C218|Anal_Canal|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C210-C212,C218|Anal_Canal|880|Sarcoma|8800/3|Sarcoma
C210-C212,C218|Anal_Canal|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C210-C212,C218|Anal_Canal|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C210-C212,C218|Anal_Canal|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C210-C212,C218|Anal_Canal|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C210-C212,C218|Anal_Canal|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C210-C212,C218|Anal_Canal|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C210-C212,C218|Anal_Canal|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C210-C212,C218|Anal_Canal|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C210-C212,C218|Anal_Canal|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C210-C212,C218|Anal_Canal|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C210-C212,C218|Anal_Canal|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C210-C212,C218|Anal_Canal|959|Lymphoma|9590/3|Lymphoma
C210-C212,C218|Anal_Canal|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C210-C212,C218|Anal_Canal|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C210-C212,C218|Anal_Canal|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C210-C212,C218|Anal_Canal|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C210-C212,C218|Anal_Canal|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C210-C212,C218|Anal_Canal|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C210-C212,C218|Anal_Canal|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C210-C212,C218|Anal_Canal|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C210-C212,C218|Anal_Canal|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C210-C212,C218|Anal_Canal|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C210-C212,C218|Anal_Canal|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C210-C212,C218|Anal_Canal|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C210-C212,C218|Anal_Canal|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C210-C212,C218|Anal_Canal|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C210-C212,C218|Anal_Canal|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C210-C212,C218|Anal_Canal|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C210-C212,C218|Anal_Canal|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C210-C212,C218|Anal_Canal|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C210-C212,C218|Anal_Canal|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C210-C212,C218|Anal_Canal|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C210-C212,C218|Anal_Canal|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C210-C212,C218|Anal_Canal|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C210-C212,C218|Anal_Canal|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C210-C212,C218|Anal_Canal|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C210-C212,C218|Anal_Canal|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C210-C212,C218|Anal_Canal|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C210-C212,C218|Anal_Canal|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C210-C212,C218|Anal_Canal|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C210-C212,C218|Anal_Canal|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C210-C212,C218|Anal_Canal|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C210-C212,C218|Anal_Canal|973|Plasmacytoma|9731/3|Plasmacytoma
C210-C212,C218|Anal_Canal|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C210-C212,C218|Anal_Canal|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C210-C212,C218|Anal_Canal|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C210-C212,C218|Anal_Canal|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C210-C212,C218|Anal_Canal|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C210-C212,C218|Anal_Canal|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C210-C212,C218|Anal_Canal|975|Neoplasm|9750/3|Malignant_Histiocytosis
C210-C212,C218|Anal_Canal|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C210-C212,C218|Anal_Canal|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C210-C212,C218|Anal_Canal|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C210-C212,C218|Anal_Canal|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C210-C212,C218|Anal_Canal|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C210-C212,C218|Anal_Canal|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C210-C212,C218|Anal_Canal|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C210-C212,C218|Anal_Canal|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C210-C212,C218|Anal_Canal|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C210-C212,C218|Anal_Canal|981|Neoplasm|9812/3|Lymphoma
C210-C212,C218|Anal_Canal|981|Neoplasm|9813/3|Lymphoma
C210-C212,C218|Anal_Canal|981|Neoplasm|9814/3|Lymphoma
C210-C212,C218|Anal_Canal|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C210-C212,C218|Anal_Canal|981|Neoplasm|9816/3|Hypodiploid_ALL
C210-C212,C218|Anal_Canal|981|Neoplasm|9817/3|Lymphoma
C210-C212,C218|Anal_Canal|981|Neoplasm|9818/3|Lymphoma
C210-C212,C218|Anal_Canal|981|Neoplasm|9819/3|Leukemia__B_Cell
C210-C212,C218|Anal_Canal|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C210-C212,C218|Anal_Canal|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C210-C212,C218|Anal_Canal|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C210-C212,C218|Anal_Canal|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C210-C212,C218|Anal_Canal|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C210-C212,C218|Anal_Canal|997|Neoplasm|9971/3|Polymorphic_PTLD
C210-C212,C218|Anal_Canal|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C220|Liver|800|Neoplasm|8000/3|Malignant_Neoplasm
C220|Liver|800|Neoplasm|8001/3|Malignant_Cell
C220|Liver|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C220|Liver|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C220|Liver|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C220|Liver|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C220|Liver|801|Carcinoma|8010/2|In_Situ_Cancer
C220|Liver|801|Carcinoma|8010/3|Carcinoma
C220|Liver|801|Carcinoma|8011/3|Malignant_Epithelioma
C220|Liver|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C220|Liver|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C220|Liver|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C220|Liver|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C220|Liver|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C220|Liver|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C220|Liver|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C220|Liver|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C220|Liver|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C220|Liver|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C220|Liver|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C220|Liver|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C220|Liver|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C220|Liver|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C220|Liver|814|Adenocarcinoma|8140/3|Adenocarcinoma
C220|Liver|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C220|Liver|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C220|Liver|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C220|Liver|816|Cholangiocarcinoma|8160/3|Cholangiocarcinoma
C220|Liver|816|Cholangiocarcinoma|8161/3|Bile_Duct_Cystadenocarcinoma
C220|Liver|817|Hepatocellular_Carcinoma|8170/3|Hepatocellular_Carcinoma
C220|Liver|817|Hepatocellular_Carcinoma|8171/3|Fibrolamellar_Carcinoma
C220|Liver|817|Hepatocellular_Carcinoma|8172/3|Scirrhous_Hepatocellular_Carcinoma
C220|Liver|817|Hepatocellular_Carcinoma|8173/3|Hepatocellular_Carcinoma
C220|Liver|817|Hepatocellular_Carcinoma|8174/3|Hepatocellular_Carcinoma
C220|Liver|817|Hepatocellular_Carcinoma|8175/3|Hepatocellular_Carcinoma
C220|Liver|818|Intrahepatic_Cholangiocarcinoma|8180/3|Cholangiocarcinoma
C220|Liver|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C220|Liver|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C220|Liver|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C220|Liver|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C220|Liver|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C220|Liver|850|Ductal_Carcinoma|8500/2|Ductal_Breast_Carcinoma_In_Situ
C220|Liver|850|Ductal_Carcinoma|8500/3|Invasive_Carcinoma
C220|Liver|850|Ductal_Carcinoma|8501/2|Comedocarcinoma
C220|Liver|850|Ductal_Carcinoma|8501/3|Comedocarcinoma
C220|Liver|850|Ductal_Carcinoma|8503/2|Intraductal_Papillary_Breast_Carcinoma
C220|Liver|850|Ductal_Carcinoma|8503/3|Intraductal_Papillary_Breast_Carcinoma
C220|Liver|850|Ductal_Carcinoma|8504/2|Intracystic_Papillary_Breast_Carcinoma
C220|Liver|850|Ductal_Carcinoma|8504/3|Intracystic_Papillary_Breast_Carcinoma
C220|Liver|850|Ductal_Carcinoma|8507/2|Micropapillary_Carcinoma
C220|Liver|850|Ductal_Carcinoma|8508/3|Carcinoma
C220|Liver|880|Sarcoma|8800/3|Sarcoma
C220|Liver|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C220|Liver|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C220|Liver|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C220|Liver|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C220|Liver|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C220|Liver|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C220|Liver|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C220|Liver|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C220|Liver|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C220|Liver|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C220|Liver|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C220|Liver|897|Hepatoblastoma|8970/3|Hepatoblastoma
C220|Liver|898|Carcinosarcoma|8980/3|Carcinosarcoma
C220|Liver|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C220|Liver|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C220|Liver|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C220|Liver|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C220|Liver|912|Neoplasms__Vascular_Tissue|9124/3|Kupffer_Cell_Sarcoma
C220|Liver|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C220|Liver|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C220|Liver|959|Lymphoma|9590/3|Lymphoma
C220|Liver|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C220|Liver|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C220|Liver|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C220|Liver|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C220|Liver|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C220|Liver|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C220|Liver|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C220|Liver|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C220|Liver|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C220|Liver|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C220|Liver|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C220|Liver|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C220|Liver|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C220|Liver|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C220|Liver|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C220|Liver|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C220|Liver|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C220|Liver|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C220|Liver|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C220|Liver|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C220|Liver|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C220|Liver|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C220|Liver|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C220|Liver|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C220|Liver|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C220|Liver|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C220|Liver|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C220|Liver|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C220|Liver|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C220|Liver|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C220|Liver|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C220|Liver|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C220|Liver|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C220|Liver|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C220|Liver|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C220|Liver|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C220|Liver|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C220|Liver|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C220|Liver|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C220|Liver|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C220|Liver|973|Plasmacytoma|9731/3|Plasmacytoma
C220|Liver|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C220|Liver|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C220|Liver|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C220|Liver|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C220|Liver|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C220|Liver|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C220|Liver|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C220|Liver|975|Neoplasm|9750/3|Malignant_Histiocytosis
C220|Liver|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C220|Liver|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C220|Liver|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C220|Liver|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C220|Liver|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C220|Liver|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C220|Liver|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C220|Liver|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C220|Liver|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C220|Liver|981|Neoplasm|9812/3|Lymphoma
C220|Liver|981|Neoplasm|9813/3|Lymphoma
C220|Liver|981|Neoplasm|9814/3|Lymphoma
C220|Liver|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C220|Liver|981|Neoplasm|9816/3|Hypodiploid_ALL
C220|Liver|981|Neoplasm|9817/3|Lymphoma
C220|Liver|981|Neoplasm|9818/3|Lymphoma
C220|Liver|981|Neoplasm|9819/3|Leukemia__B_Cell
C220|Liver|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C220|Liver|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C220|Liver|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C220|Liver|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C220|Liver|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C220|Liver|997|Neoplasm|9971/3|Polymorphic_PTLD
C220|Liver|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C221|Intrahepatic_Bile_Duct|800|Neoplasm|8000/3|Malignant_Neoplasm
C221|Intrahepatic_Bile_Duct|800|Neoplasm|8001/3|Malignant_Cell
C221|Intrahepatic_Bile_Duct|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C221|Intrahepatic_Bile_Duct|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C221|Intrahepatic_Bile_Duct|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C221|Intrahepatic_Bile_Duct|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C221|Intrahepatic_Bile_Duct|801|Carcinoma|8010/2|In_Situ_Cancer
C221|Intrahepatic_Bile_Duct|801|Carcinoma|8010/3|Carcinoma
C221|Intrahepatic_Bile_Duct|801|Carcinoma|8011/3|Malignant_Epithelioma
C221|Intrahepatic_Bile_Duct|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C221|Intrahepatic_Bile_Duct|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C221|Intrahepatic_Bile_Duct|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C221|Intrahepatic_Bile_Duct|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C221|Intrahepatic_Bile_Duct|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C221|Intrahepatic_Bile_Duct|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C221|Intrahepatic_Bile_Duct|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C221|Intrahepatic_Bile_Duct|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C221|Intrahepatic_Bile_Duct|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C221|Intrahepatic_Bile_Duct|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C221|Intrahepatic_Bile_Duct|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C221|Intrahepatic_Bile_Duct|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C221|Intrahepatic_Bile_Duct|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C221|Intrahepatic_Bile_Duct|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C221|Intrahepatic_Bile_Duct|814|Adenocarcinoma|8140/3|Adenocarcinoma
C221|Intrahepatic_Bile_Duct|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C221|Intrahepatic_Bile_Duct|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C221|Intrahepatic_Bile_Duct|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C221|Intrahepatic_Bile_Duct|816|Cholangiocarcinoma|8160/3|Cholangiocarcinoma
C221|Intrahepatic_Bile_Duct|816|Cholangiocarcinoma|8161/3|Bile_Duct_Cystadenocarcinoma
C221|Intrahepatic_Bile_Duct|816|Cholangiocarcinoma|8162/3|Hilar_Cholangiocarcinoma
C221|Intrahepatic_Bile_Duct|817|Hepatocellular_Carcinoma|8170/3|Hepatocellular_Carcinoma
C221|Intrahepatic_Bile_Duct|817|Hepatocellular_Carcinoma|8171/3|Fibrolamellar_Carcinoma
C221|Intrahepatic_Bile_Duct|817|Hepatocellular_Carcinoma|8172/3|Scirrhous_Hepatocellular_Carcinoma
C221|Intrahepatic_Bile_Duct|817|Hepatocellular_Carcinoma|8173/3|Hepatocellular_Carcinoma
C221|Intrahepatic_Bile_Duct|817|Hepatocellular_Carcinoma|8174/3|Hepatocellular_Carcinoma
C221|Intrahepatic_Bile_Duct|817|Hepatocellular_Carcinoma|8175/3|Hepatocellular_Carcinoma
C221|Intrahepatic_Bile_Duct|818|Intrahepatic_Cholangiocarcinoma|8180/3|Cholangiocarcinoma
C221|Intrahepatic_Bile_Duct|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C221|Intrahepatic_Bile_Duct|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C221|Intrahepatic_Bile_Duct|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C221|Intrahepatic_Bile_Duct|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C221|Intrahepatic_Bile_Duct|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8500/2|Ductal_Breast_Carcinoma_In_Situ
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8500/3|Invasive_Carcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8501/2|Comedocarcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8501/3|Comedocarcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8503/2|Intraductal_Papillary_Breast_Carcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8503/3|Intraductal_Papillary_Breast_Carcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8504/2|Intracystic_Papillary_Breast_Carcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8504/3|Intracystic_Papillary_Breast_Carcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8507/2|Micropapillary_Carcinoma
C221|Intrahepatic_Bile_Duct|850|Ductal_Carcinoma|8508/3|Carcinoma
C221|Intrahepatic_Bile_Duct|880|Sarcoma|8800/3|Sarcoma
C221|Intrahepatic_Bile_Duct|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C221|Intrahepatic_Bile_Duct|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C221|Intrahepatic_Bile_Duct|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C221|Intrahepatic_Bile_Duct|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C221|Intrahepatic_Bile_Duct|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C221|Intrahepatic_Bile_Duct|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C221|Intrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C221|Intrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C221|Intrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C221|Intrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C221|Intrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C221|Intrahepatic_Bile_Duct|898|Carcinosarcoma|8980/3|Carcinosarcoma
C221|Intrahepatic_Bile_Duct|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C221|Intrahepatic_Bile_Duct|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C221|Intrahepatic_Bile_Duct|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C221|Intrahepatic_Bile_Duct|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C221|Intrahepatic_Bile_Duct|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C221|Intrahepatic_Bile_Duct|959|Lymphoma|9590/3|Lymphoma
C221|Intrahepatic_Bile_Duct|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C221|Intrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C221|Intrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C221|Intrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C221|Intrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C221|Intrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C221|Intrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C221|Intrahepatic_Bile_Duct|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C221|Intrahepatic_Bile_Duct|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C221|Intrahepatic_Bile_Duct|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C221|Intrahepatic_Bile_Duct|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C221|Intrahepatic_Bile_Duct|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C221|Intrahepatic_Bile_Duct|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C221|Intrahepatic_Bile_Duct|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C221|Intrahepatic_Bile_Duct|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C221|Intrahepatic_Bile_Duct|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C221|Intrahepatic_Bile_Duct|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C221|Intrahepatic_Bile_Duct|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C221|Intrahepatic_Bile_Duct|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C221|Intrahepatic_Bile_Duct|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C221|Intrahepatic_Bile_Duct|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C221|Intrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C221|Intrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C221|Intrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C221|Intrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C221|Intrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C221|Intrahepatic_Bile_Duct|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C221|Intrahepatic_Bile_Duct|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C221|Intrahepatic_Bile_Duct|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C221|Intrahepatic_Bile_Duct|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C221|Intrahepatic_Bile_Duct|973|Plasmacytoma|9731/3|Plasmacytoma
C221|Intrahepatic_Bile_Duct|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C221|Intrahepatic_Bile_Duct|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C221|Intrahepatic_Bile_Duct|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C221|Intrahepatic_Bile_Duct|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C221|Intrahepatic_Bile_Duct|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C221|Intrahepatic_Bile_Duct|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C221|Intrahepatic_Bile_Duct|975|Neoplasm|9750/3|Malignant_Histiocytosis
C221|Intrahepatic_Bile_Duct|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C221|Intrahepatic_Bile_Duct|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C221|Intrahepatic_Bile_Duct|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C221|Intrahepatic_Bile_Duct|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C221|Intrahepatic_Bile_Duct|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C221|Intrahepatic_Bile_Duct|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C221|Intrahepatic_Bile_Duct|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C221|Intrahepatic_Bile_Duct|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9812/3|Lymphoma
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9813/3|Lymphoma
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9814/3|Lymphoma
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9816/3|Hypodiploid_ALL
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9817/3|Lymphoma
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9818/3|Lymphoma
C221|Intrahepatic_Bile_Duct|981|Neoplasm|9819/3|Leukemia__B_Cell
C221|Intrahepatic_Bile_Duct|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C221|Intrahepatic_Bile_Duct|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C221|Intrahepatic_Bile_Duct|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C221|Intrahepatic_Bile_Duct|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C221|Intrahepatic_Bile_Duct|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C221|Intrahepatic_Bile_Duct|997|Neoplasm|9971/3|Polymorphic_PTLD
C221|Intrahepatic_Bile_Duct|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C239-C241,C248-C249|Extrahepatic_Bile_Duct|800|Neoplasm|8000/3|Malignant_Neoplasm
C239-C241,C248-C249|Extrahepatic_Bile_Duct|800|Neoplasm|8001/3|Malignant_Cell
C239-C241,C248-C249|Extrahepatic_Bile_Duct|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C239-C241,C248-C249|Extrahepatic_Bile_Duct|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C239-C241,C248-C249|Extrahepatic_Bile_Duct|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C239-C241,C248-C249|Extrahepatic_Bile_Duct|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C239-C241,C248-C249|Extrahepatic_Bile_Duct|801|Carcinoma|8010/2|In_Situ_Cancer
C239-C241,C248-C249|Extrahepatic_Bile_Duct|801|Carcinoma|8010/3|Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|801|Carcinoma|8011/3|Malignant_Epithelioma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C239-C241,C248-C249|Extrahepatic_Bile_Duct|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C239-C241,C248-C249|Extrahepatic_Bile_Duct|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C239-C241,C248-C249|Extrahepatic_Bile_Duct|814|Adenocarcinoma|8140/3|Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C239-C241,C248-C249|Extrahepatic_Bile_Duct|816|Cholangiocarcinoma|8160/3|Cholangiocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|816|Cholangiocarcinoma|8161/3|Bile_Duct_Cystadenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|816|Cholangiocarcinoma|8162/3|Hilar_Cholangiocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|816|Cholangiocarcinoma|8163/3|Pancreatobiliary_type_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C239-C241,C248-C249|Extrahepatic_Bile_Duct|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C239-C241,C248-C249|Extrahepatic_Bile_Duct|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C239-C241,C248-C249|Extrahepatic_Bile_Duct|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8500/2|Ductal_Breast_Carcinoma_In_Situ
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8500/3|Invasive_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8501/2|Comedocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8501/3|Comedocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8503/2|Intraductal_Papillary_Breast_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8503/3|Intraductal_Papillary_Breast_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8504/2|Intracystic_Papillary_Breast_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8504/3|Intracystic_Papillary_Breast_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8507/2|Micropapillary_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|850|Ductal_Carcinoma|8508/3|Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C239-C241,C248-C249|Extrahepatic_Bile_Duct|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C239-C241,C248-C249|Extrahepatic_Bile_Duct|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|880|Sarcoma|8800/3|Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C239-C241,C248-C249|Extrahepatic_Bile_Duct|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C239-C241,C248-C249|Extrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|898|Carcinosarcoma|8980/3|Carcinosarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C239-C241,C248-C249|Extrahepatic_Bile_Duct|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|959|Lymphoma|9590/3|Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C239-C241,C248-C249|Extrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C239-C241,C248-C249|Extrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C239-C241,C248-C249|Extrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C239-C241,C248-C249|Extrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C239-C241,C248-C249|Extrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C239-C241,C248-C249|Extrahepatic_Bile_Duct|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C239-C241,C248-C249|Extrahepatic_Bile_Duct|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C239-C241,C248-C249|Extrahepatic_Bile_Duct|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C239-C241,C248-C249|Extrahepatic_Bile_Duct|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C239-C241,C248-C249|Extrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C239-C241,C248-C249|Extrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C239-C241,C248-C249|Extrahepatic_Bile_Duct|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|973|Plasmacytoma|9731/3|Plasmacytoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C239-C241,C248-C249|Extrahepatic_Bile_Duct|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C239-C241,C248-C249|Extrahepatic_Bile_Duct|975|Neoplasm|9750/3|Malignant_Histiocytosis
C239-C241,C248-C249|Extrahepatic_Bile_Duct|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C239-C241,C248-C249|Extrahepatic_Bile_Duct|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C239-C241,C248-C249|Extrahepatic_Bile_Duct|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C239-C241,C248-C249|Extrahepatic_Bile_Duct|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9812/3|Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9813/3|Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9814/3|Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9816/3|Hypodiploid_ALL
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9817/3|Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9818/3|Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|981|Neoplasm|9819/3|Leukemia__B_Cell
C239-C241,C248-C249|Extrahepatic_Bile_Duct|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C239-C241,C248-C249|Extrahepatic_Bile_Duct|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C239-C241,C248-C249|Extrahepatic_Bile_Duct|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C239-C241,C248-C249|Extrahepatic_Bile_Duct|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C239-C241,C248-C249|Extrahepatic_Bile_Duct|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C239-C241,C248-C249|Extrahepatic_Bile_Duct|997|Neoplasm|9971/3|Polymorphic_PTLD
C239-C241,C248-C249|Extrahepatic_Bile_Duct|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C250-C254,C257-C259|Pancreas|800|Neoplasm|8000/3|Malignant_Neoplasm
C250-C254,C257-C259|Pancreas|800|Neoplasm|8001/3|Malignant_Cell
C250-C254,C257-C259|Pancreas|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C250-C254,C257-C259|Pancreas|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C250-C254,C257-C259|Pancreas|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C250-C254,C257-C259|Pancreas|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C250-C254,C257-C259|Pancreas|801|Carcinoma|8010/2|In_Situ_Cancer
C250-C254,C257-C259|Pancreas|801|Carcinoma|8010/3|Carcinoma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8011/3|Malignant_Epithelioma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C250-C254,C257-C259|Pancreas|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C250-C254,C257-C259|Pancreas|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C250-C254,C257-C259|Pancreas|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C250-C254,C257-C259|Pancreas|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C250-C254,C257-C259|Pancreas|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C250-C254,C257-C259|Pancreas|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C250-C254,C257-C259|Pancreas|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C250-C254,C257-C259|Pancreas|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C250-C254,C257-C259|Pancreas|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C250-C254,C257-C259|Pancreas|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C250-C254,C257-C259|Pancreas|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8140/3|Adenocarcinoma
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C250-C254,C257-C259|Pancreas|814|Adenocarcinoma|8148/2|Intraepithelial_Neoplasia
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8150/3|Pancreatic_Endocrine_Carcinoma
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8151/3|Malignant_Pancreatic_Insulinoma
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8152/3|Malignant_Pancreatic_Glucagonoma
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8153/3|Malignant_Gastrinoma
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8154/3|Adenocarcinoma
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8155/3|Malignant_Vipoma
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8156/3|Malignant_Somatostatinoma
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8157/3|Malignant_Enteroglucagonoma
C250-C254,C257-C259|Pancreas|815|Endocrine_Gland_Neoplasms|8158/3|Neoplasm
C250-C254,C257-C259|Pancreas|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C250-C254,C257-C259|Pancreas|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C250-C254,C257-C259|Pancreas|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C250-C254,C257-C259|Pancreas|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C250-C254,C257-C259|Pancreas|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C250-C254,C257-C259|Pancreas|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C250-C254,C257-C259|Pancreas|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C250-C254,C257-C259|Pancreas|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C250-C254,C257-C259|Pancreas|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C250-C254,C257-C259|Pancreas|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C250-C254,C257-C259|Pancreas|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C250-C254,C257-C259|Pancreas|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C250-C254,C257-C259|Pancreas|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C250-C254,C257-C259|Pancreas|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C250-C254,C257-C259|Pancreas|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C250-C254,C257-C259|Pancreas|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C250-C254,C257-C259|Pancreas|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C250-C254,C257-C259|Pancreas|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C250-C254,C257-C259|Pancreas|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C250-C254,C257-C259|Pancreas|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C250-C254,C257-C259|Pancreas|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C250-C254,C257-C259|Pancreas|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C250-C254,C257-C259|Pancreas|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C250-C254,C257-C259|Pancreas|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C250-C254,C257-C259|Pancreas|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C250-C254,C257-C259|Pancreas|845|Papillary_Cystadenocarcinoma|8450/3|Papillary_Cystadenocarcinoma
C250-C254,C257-C259|Pancreas|845|Papillary_Cystadenocarcinoma|8452/3|Carcinoma
C250-C254,C257-C259|Pancreas|845|Papillary_Cystadenocarcinoma|8453/2|Mucinous_Adenocarcinoma
C250-C254,C257-C259|Pancreas|845|Papillary_Cystadenocarcinoma|8453/3|Mucinous_Adenocarcinoma
C250-C254,C257-C259|Pancreas|847|Mucinous_Cystadenocarcinoma|8470/2|Mucinous_Cystadenocarcinoma
C250-C254,C257-C259|Pancreas|847|Mucinous_Cystadenocarcinoma|8470/3|Mucinous_Cystadenocarcinoma
C250-C254,C257-C259|Pancreas|847|Mucinous_Cystadenocarcinoma|8471/3|Papillary_Mucinous_Cystadenocarcinoma
C250-C254,C257-C259|Pancreas|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C250-C254,C257-C259|Pancreas|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C250-C254,C257-C259|Pancreas|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8500/2|Ductal_Breast_Carcinoma_In_Situ
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8500/3|Invasive_Carcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8501/2|Comedocarcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8501/3|Comedocarcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8503/2|Intraductal_Papillary_Breast_Carcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8503/3|Intraductal_Papillary_Breast_Carcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8504/2|Intracystic_Papillary_Breast_Carcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8504/3|Intracystic_Papillary_Breast_Carcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8507/2|Micropapillary_Carcinoma
C250-C254,C257-C259|Pancreas|850|Ductal_Carcinoma|8508/3|Carcinoma
C250-C254,C257-C259|Pancreas|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C250-C254,C257-C259|Pancreas|851|Medullary_Carcinoma|8514/3|Ductal_Carcinoma
C250-C254,C257-C259|Pancreas|852|Intraductal_And_Lobular_Carcinoma|8521/3|Invasive_Ductal_Breast_Carcinoma
C250-C254,C257-C259|Pancreas|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C250-C254,C257-C259|Pancreas|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C250-C254,C257-C259|Pancreas|855|Acinar_Cell_Carcinoma|8552/3|Ductal_Carcinoma
C250-C254,C257-C259|Pancreas|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C250-C254,C257-C259|Pancreas|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C250-C254,C257-C259|Pancreas|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C250-C254,C257-C259|Pancreas|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C250-C254,C257-C259|Pancreas|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C250-C254,C257-C259|Pancreas|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C250-C254,C257-C259|Pancreas|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C250-C254,C257-C259|Pancreas|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C250-C254,C257-C259|Pancreas|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8800/3|Sarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C250-C254,C257-C259|Pancreas|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C250-C254,C257-C259|Pancreas|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C250-C254,C257-C259|Pancreas|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C250-C254,C257-C259|Pancreas|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C250-C254,C257-C259|Pancreas|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C250-C254,C257-C259|Pancreas|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C250-C254,C257-C259|Pancreas|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C250-C254,C257-C259|Pancreas|897|Pancreatoblastoma|8971/3|Pancreatoblastoma
C250-C254,C257-C259|Pancreas|898|Carcinosarcoma|8980/3|Carcinosarcoma
C250-C254,C257-C259|Pancreas|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C250-C254,C257-C259|Pancreas|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C250-C254,C257-C259|Pancreas|959|Lymphoma|9590/3|Lymphoma
C250-C254,C257-C259|Pancreas|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C250-C254,C257-C259|Pancreas|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C250-C254,C257-C259|Pancreas|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C250-C254,C257-C259|Pancreas|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C250-C254,C257-C259|Pancreas|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C250-C254,C257-C259|Pancreas|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C250-C254,C257-C259|Pancreas|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C250-C254,C257-C259|Pancreas|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C250-C254,C257-C259|Pancreas|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C250-C254,C257-C259|Pancreas|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C250-C254,C257-C259|Pancreas|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C250-C254,C257-C259|Pancreas|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C250-C254,C257-C259|Pancreas|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C250-C254,C257-C259|Pancreas|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C250-C254,C257-C259|Pancreas|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C250-C254,C257-C259|Pancreas|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C250-C254,C257-C259|Pancreas|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C250-C254,C257-C259|Pancreas|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C250-C254,C257-C259|Pancreas|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C250-C254,C257-C259|Pancreas|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C250-C254,C257-C259|Pancreas|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C250-C254,C257-C259|Pancreas|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C250-C254,C257-C259|Pancreas|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C250-C254,C257-C259|Pancreas|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C250-C254,C257-C259|Pancreas|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C250-C254,C257-C259|Pancreas|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C250-C254,C257-C259|Pancreas|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C250-C254,C257-C259|Pancreas|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C250-C254,C257-C259|Pancreas|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9731/3|Plasmacytoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C250-C254,C257-C259|Pancreas|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C250-C254,C257-C259|Pancreas|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C250-C254,C257-C259|Pancreas|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C250-C254,C257-C259|Pancreas|975|Neoplasm|9750/3|Malignant_Histiocytosis
C250-C254,C257-C259|Pancreas|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C250-C254,C257-C259|Pancreas|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C250-C254,C257-C259|Pancreas|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C250-C254,C257-C259|Pancreas|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C250-C254,C257-C259|Pancreas|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C250-C254,C257-C259|Pancreas|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C250-C254,C257-C259|Pancreas|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C250-C254,C257-C259|Pancreas|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C250-C254,C257-C259|Pancreas|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C250-C254,C257-C259|Pancreas|981|Neoplasm|9812/3|Lymphoma
C250-C254,C257-C259|Pancreas|981|Neoplasm|9813/3|Lymphoma
C250-C254,C257-C259|Pancreas|981|Neoplasm|9814/3|Lymphoma
C250-C254,C257-C259|Pancreas|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C250-C254,C257-C259|Pancreas|981|Neoplasm|9816/3|Hypodiploid_ALL
C250-C254,C257-C259|Pancreas|981|Neoplasm|9817/3|Lymphoma
C250-C254,C257-C259|Pancreas|981|Neoplasm|9818/3|Lymphoma
C250-C254,C257-C259|Pancreas|981|Neoplasm|9819/3|Leukemia__B_Cell
C250-C254,C257-C259|Pancreas|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C250-C254,C257-C259|Pancreas|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C250-C254,C257-C259|Pancreas|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C250-C254,C257-C259|Pancreas|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C250-C254,C257-C259|Pancreas|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C250-C254,C257-C259|Pancreas|997|Neoplasm|9971/3|Polymorphic_PTLD
C250-C254,C257-C259|Pancreas|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C260,C268-C269|Entire_Digestive_Organ|800|Neoplasm|8000/3|Malignant_Neoplasm
C260,C268-C269|Entire_Digestive_Organ|800|Neoplasm|8001/3|Malignant_Cell
C260,C268-C269|Entire_Digestive_Organ|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C260,C268-C269|Entire_Digestive_Organ|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C260,C268-C269|Entire_Digestive_Organ|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C260,C268-C269|Entire_Digestive_Organ|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C260,C268-C269|Entire_Digestive_Organ|801|Carcinoma|8010/2|In_Situ_Cancer
C260,C268-C269|Entire_Digestive_Organ|801|Carcinoma|8010/3|Carcinoma
C260,C268-C269|Entire_Digestive_Organ|801|Carcinoma|8011/3|Malignant_Epithelioma
C260,C268-C269|Entire_Digestive_Organ|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C260,C268-C269|Entire_Digestive_Organ|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C260,C268-C269|Entire_Digestive_Organ|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C260,C268-C269|Entire_Digestive_Organ|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C260,C268-C269|Entire_Digestive_Organ|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|813|Carcinoma|8130/2|Carcinoma
C260,C268-C269|Entire_Digestive_Organ|813|Carcinoma|8130/3|Carcinoma
C260,C268-C269|Entire_Digestive_Organ|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C260,C268-C269|Entire_Digestive_Organ|814|Adenocarcinoma|8140/3|Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C260,C268-C269|Entire_Digestive_Organ|815|Endocrine_Gland_Neoplasms|8152/3|Malignant_Pancreatic_Glucagonoma
C260,C268-C269|Entire_Digestive_Organ|815|Endocrine_Gland_Neoplasms|8153/3|Malignant_Gastrinoma
C260,C268-C269|Entire_Digestive_Organ|815|Endocrine_Gland_Neoplasms|8156/3|Malignant_Somatostatinoma
C260,C268-C269|Entire_Digestive_Organ|815|Endocrine_Gland_Neoplasms|8157/3|Malignant_Enteroglucagonoma
C260,C268-C269|Entire_Digestive_Organ|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C260,C268-C269|Entire_Digestive_Organ|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C260,C268-C269|Entire_Digestive_Organ|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C260,C268-C269|Entire_Digestive_Organ|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C260,C268-C269|Entire_Digestive_Organ|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C260,C268-C269|Entire_Digestive_Organ|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C260,C268-C269|Entire_Digestive_Organ|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C260,C268-C269|Entire_Digestive_Organ|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C260,C268-C269|Entire_Digestive_Organ|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C260,C268-C269|Entire_Digestive_Organ|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C260,C268-C269|Entire_Digestive_Organ|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C260,C268-C269|Entire_Digestive_Organ|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C260,C268-C269|Entire_Digestive_Organ|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C260,C268-C269|Entire_Digestive_Organ|825|Bronchioloalveolar_Adenocarcinoma|8251/3|Bronchioloalveolar_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C260,C268-C269|Entire_Digestive_Organ|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C260,C268-C269|Entire_Digestive_Organ|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C260,C268-C269|Entire_Digestive_Organ|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C260,C268-C269|Entire_Digestive_Organ|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C260,C268-C269|Entire_Digestive_Organ|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C260,C268-C269|Entire_Digestive_Organ|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|850|Ductal_Carcinoma|8503/2|Intraductal_Papillary_Breast_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|850|Ductal_Carcinoma|8503/3|Intraductal_Papillary_Breast_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|850|Ductal_Carcinoma|8504/2|Intracystic_Papillary_Breast_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|850|Ductal_Carcinoma|8504/3|Intracystic_Papillary_Breast_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|852|Intraductal_And_Lobular_Carcinoma|8521/3|Invasive_Ductal_Breast_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C260,C268-C269|Entire_Digestive_Organ|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C260,C268-C269|Entire_Digestive_Organ|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C260,C268-C269|Entire_Digestive_Organ|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C260,C268-C269|Entire_Digestive_Organ|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C260,C268-C269|Entire_Digestive_Organ|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C260,C268-C269|Entire_Digestive_Organ|872|Melanoma|8720/3|Melanoma
C260,C268-C269|Entire_Digestive_Organ|872|Melanoma|8721/3|Nodular_Melanoma
C260,C268-C269|Entire_Digestive_Organ|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C260,C268-C269|Entire_Digestive_Organ|872|Melanoma|8723/3|Regressing_Melanoma
C260,C268-C269|Entire_Digestive_Organ|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C260,C268-C269|Entire_Digestive_Organ|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C260,C268-C269|Entire_Digestive_Organ|874|Nevus|8745/3|Desmoplastic_Melanoma
C260,C268-C269|Entire_Digestive_Organ|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C260,C268-C269|Entire_Digestive_Organ|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C260,C268-C269|Entire_Digestive_Organ|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C260,C268-C269|Entire_Digestive_Organ|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C260,C268-C269|Entire_Digestive_Organ|880|Sarcoma|8800/3|Sarcoma
C260,C268-C269|Entire_Digestive_Organ|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C260,C268-C269|Entire_Digestive_Organ|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C260,C268-C269|Entire_Digestive_Organ|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C260,C268-C269|Entire_Digestive_Organ|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C260,C268-C269|Entire_Digestive_Organ|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C260,C268-C269|Entire_Digestive_Organ|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C260,C268-C269|Entire_Digestive_Organ|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C260,C268-C269|Entire_Digestive_Organ|882|Sarcoma|8825/3|Sarcoma
C260,C268-C269|Entire_Digestive_Organ|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C260,C268-C269|Entire_Digestive_Organ|884|Myxosarcoma|8840/3|Myxosarcoma
C260,C268-C269|Entire_Digestive_Organ|885|Liposarcoma|8850/3|Liposarcoma
C260,C268-C269|Entire_Digestive_Organ|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C260,C268-C269|Entire_Digestive_Organ|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C260,C268-C269|Entire_Digestive_Organ|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C260,C268-C269|Entire_Digestive_Organ|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C260,C268-C269|Entire_Digestive_Organ|885|Liposarcoma|8855/3|Liposarcoma
C260,C268-C269|Entire_Digestive_Organ|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C260,C268-C269|Entire_Digestive_Organ|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C260,C268-C269|Entire_Digestive_Organ|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C260,C268-C269|Entire_Digestive_Organ|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C260,C268-C269|Entire_Digestive_Organ|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|893|Stromal_Sarcoma|8936/3|High_Risk_Gastrointestinal_Stromal_Tumor
C260,C268-C269|Entire_Digestive_Organ|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C260,C268-C269|Entire_Digestive_Organ|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C260,C268-C269|Entire_Digestive_Organ|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C260,C268-C269|Entire_Digestive_Organ|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C260,C268-C269|Entire_Digestive_Organ|898|Carcinosarcoma|8980/3|Carcinosarcoma
C260,C268-C269|Entire_Digestive_Organ|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C260,C268-C269|Entire_Digestive_Organ|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C260,C268-C269|Entire_Digestive_Organ|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C260,C268-C269|Entire_Digestive_Organ|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C260,C268-C269|Entire_Digestive_Organ|904|Synovial_Sarcoma|9040/3|Synovial_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|904|Synovial_Sarcoma|9041/3|Spindle_Cell_Synovial_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|904|Synovial_Sarcoma|9042/3|Epithelial_Synovial_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|904|Synovial_Sarcoma|9043/3|Biphasic_Synovial_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|904|Synovial_Sarcoma|9044/3|Clear_Cell_Sarcoma_Of_Soft_Tissue_C0206651
C260,C268-C269|Entire_Digestive_Organ|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C260,C268-C269|Entire_Digestive_Organ|906|Germ_Cell_Tumor|9064/3|Germinoma
C260,C268-C269|Entire_Digestive_Organ|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C260,C268-C269|Entire_Digestive_Organ|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C260,C268-C269|Entire_Digestive_Organ|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C260,C268-C269|Entire_Digestive_Organ|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C260,C268-C269|Entire_Digestive_Organ|908|Teratoma|9080/3|Immature_Teratoma
C260,C268-C269|Entire_Digestive_Organ|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C260,C268-C269|Entire_Digestive_Organ|908|Teratoma|9082/3|Immature_Teratoma
C260,C268-C269|Entire_Digestive_Organ|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C260,C268-C269|Entire_Digestive_Organ|908|Teratoma|9084/3|Teratoma
C260,C268-C269|Entire_Digestive_Organ|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C260,C268-C269|Entire_Digestive_Organ|910|Choriocarcinoma|9100/3|Choriocarcinoma
C260,C268-C269|Entire_Digestive_Organ|910|Choriocarcinoma|9101/3|Choriocarcinoma
C260,C268-C269|Entire_Digestive_Organ|910|Choriocarcinoma|9105/3|Epithelioid_Trophoblastic_Tumor
C260,C268-C269|Entire_Digestive_Organ|911|Mesonephroma|9110/3|Mesonephroma
C260,C268-C269|Entire_Digestive_Organ|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C260,C268-C269|Entire_Digestive_Organ|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C260,C268-C269|Entire_Digestive_Organ|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C260,C268-C269|Entire_Digestive_Organ|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C260,C268-C269|Entire_Digestive_Organ|917|Lymphangiosarcoma|9170/3|Lymphangiosarcoma
C260,C268-C269|Entire_Digestive_Organ|925|Bone_Neoplasm|9251/3|Giant_Cell_Tumor_Of_Soft_Tissue
C260,C268-C269|Entire_Digestive_Organ|925|Bone_Neoplasm|9252/3|Malignant_Tenosynovial_Giant_Cell_Tumor
C260,C268-C269|Entire_Digestive_Organ|937|Chordoma|9370/3|Chordoma
C260,C268-C269|Entire_Digestive_Organ|937|Chordoma|9371/3|Chondroid_Chordoma
C260,C268-C269|Entire_Digestive_Organ|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C260,C268-C269|Entire_Digestive_Organ|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C260,C268-C269|Entire_Digestive_Organ|950|Neuroblastoma|9500/3|Neuroblastoma
C260,C268-C269|Entire_Digestive_Organ|950|Neuroblastoma|9501/3|Medulloepithelioma
C260,C268-C269|Entire_Digestive_Organ|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C260,C268-C269|Entire_Digestive_Organ|950|Neuroblastoma|9503/3|Neuroepithelioma
C260,C268-C269|Entire_Digestive_Organ|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C260,C268-C269|Entire_Digestive_Organ|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C260,C268-C269|Entire_Digestive_Organ|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C260,C268-C269|Entire_Digestive_Organ|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C260,C268-C269|Entire_Digestive_Organ|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C260,C268-C269|Entire_Digestive_Organ|957|Perineurioma|9571/3|Malignant_Perineurioma
C260,C268-C269|Entire_Digestive_Organ|959|Lymphoma|9590/3|Lymphoma
C260,C268-C269|Entire_Digestive_Organ|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C260,C268-C269|Entire_Digestive_Organ|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C260,C268-C269|Entire_Digestive_Organ|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C260,C268-C269|Entire_Digestive_Organ|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C260,C268-C269|Entire_Digestive_Organ|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C260,C268-C269|Entire_Digestive_Organ|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C260,C268-C269|Entire_Digestive_Organ|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C260,C268-C269|Entire_Digestive_Organ|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C260,C268-C269|Entire_Digestive_Organ|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C260,C268-C269|Entire_Digestive_Organ|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C260,C268-C269|Entire_Digestive_Organ|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C260,C268-C269|Entire_Digestive_Organ|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C260,C268-C269|Entire_Digestive_Organ|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C260,C268-C269|Entire_Digestive_Organ|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C260,C268-C269|Entire_Digestive_Organ|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C260,C268-C269|Entire_Digestive_Organ|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|973|Plasmacytoma|9731/3|Plasmacytoma
C260,C268-C269|Entire_Digestive_Organ|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C260,C268-C269|Entire_Digestive_Organ|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C260,C268-C269|Entire_Digestive_Organ|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C260,C268-C269|Entire_Digestive_Organ|975|Neoplasm|9750/3|Malignant_Histiocytosis
C260,C268-C269|Entire_Digestive_Organ|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C260,C268-C269|Entire_Digestive_Organ|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C260,C268-C269|Entire_Digestive_Organ|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C260,C268-C269|Entire_Digestive_Organ|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C260,C268-C269|Entire_Digestive_Organ|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9812/3|Lymphoma
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9813/3|Lymphoma
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9814/3|Lymphoma
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9816/3|Hypodiploid_ALL
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9817/3|Lymphoma
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9818/3|Lymphoma
C260,C268-C269|Entire_Digestive_Organ|981|Neoplasm|9819/3|Leukemia__B_Cell
C260,C268-C269|Entire_Digestive_Organ|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C260,C268-C269|Entire_Digestive_Organ|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C260,C268-C269|Entire_Digestive_Organ|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C260,C268-C269|Entire_Digestive_Organ|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C260,C268-C269|Entire_Digestive_Organ|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C260,C268-C269|Entire_Digestive_Organ|997|Neoplasm|9971/3|Polymorphic_PTLD
C260,C268-C269|Entire_Digestive_Organ|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C300|Nasal_Cartilage|800|Neoplasm|8000/3|Malignant_Neoplasm
C300|Nasal_Cartilage|800|Neoplasm|8001/3|Malignant_Cell
C300|Nasal_Cartilage|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C300|Nasal_Cartilage|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C300|Nasal_Cartilage|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C300|Nasal_Cartilage|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C300|Nasal_Cartilage|801|Carcinoma|8010/2|In_Situ_Cancer
C300|Nasal_Cartilage|801|Carcinoma|8010/3|Carcinoma
C300|Nasal_Cartilage|801|Carcinoma|8011/3|Malignant_Epithelioma
C300|Nasal_Cartilage|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C300|Nasal_Cartilage|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C300|Nasal_Cartilage|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C300|Nasal_Cartilage|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C300|Nasal_Cartilage|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C300|Nasal_Cartilage|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C300|Nasal_Cartilage|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C300|Nasal_Cartilage|802|Carcinoma|8023/3|NUT_Carcinoma
C300|Nasal_Cartilage|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C300|Nasal_Cartilage|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C300|Nasal_Cartilage|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C300|Nasal_Cartilage|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C300|Nasal_Cartilage|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C300|Nasal_Cartilage|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C300|Nasal_Cartilage|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C300|Nasal_Cartilage|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C300|Nasal_Cartilage|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C300|Nasal_Cartilage|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C300|Nasal_Cartilage|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C300|Nasal_Cartilage|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C300|Nasal_Cartilage|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C300|Nasal_Cartilage|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C300|Nasal_Cartilage|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C300|Nasal_Cartilage|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C300|Nasal_Cartilage|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C300|Nasal_Cartilage|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C300|Nasal_Cartilage|813|Carcinoma|8130/2|Carcinoma
C300|Nasal_Cartilage|813|Carcinoma|8130/3|Carcinoma
C300|Nasal_Cartilage|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C300|Nasal_Cartilage|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C300|Nasal_Cartilage|814|Adenocarcinoma|8140/3|Adenocarcinoma
C300|Nasal_Cartilage|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C300|Nasal_Cartilage|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C300|Nasal_Cartilage|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C300|Nasal_Cartilage|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C300|Nasal_Cartilage|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C300|Nasal_Cartilage|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C300|Nasal_Cartilage|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C300|Nasal_Cartilage|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C300|Nasal_Cartilage|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C300|Nasal_Cartilage|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C300|Nasal_Cartilage|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C300|Nasal_Cartilage|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C300|Nasal_Cartilage|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C300|Nasal_Cartilage|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C300|Nasal_Cartilage|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C300|Nasal_Cartilage|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C300|Nasal_Cartilage|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C300|Nasal_Cartilage|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C300|Nasal_Cartilage|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C300|Nasal_Cartilage|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C300|Nasal_Cartilage|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C300|Nasal_Cartilage|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C300|Nasal_Cartilage|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C300|Nasal_Cartilage|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C300|Nasal_Cartilage|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C300|Nasal_Cartilage|872|Melanoma|8720/3|Melanoma
C300|Nasal_Cartilage|872|Melanoma|8721/3|Nodular_Melanoma
C300|Nasal_Cartilage|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C300|Nasal_Cartilage|872|Melanoma|8723/3|Regressing_Melanoma
C300|Nasal_Cartilage|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C300|Nasal_Cartilage|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C300|Nasal_Cartilage|874|Nevus|8745/3|Desmoplastic_Melanoma
C300|Nasal_Cartilage|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C300|Nasal_Cartilage|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C300|Nasal_Cartilage|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C300|Nasal_Cartilage|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C300|Nasal_Cartilage|880|Sarcoma|8800/3|Sarcoma
C300|Nasal_Cartilage|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C300|Nasal_Cartilage|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C300|Nasal_Cartilage|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C300|Nasal_Cartilage|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C300|Nasal_Cartilage|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C300|Nasal_Cartilage|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C300|Nasal_Cartilage|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C300|Nasal_Cartilage|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C300|Nasal_Cartilage|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C300|Nasal_Cartilage|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C300|Nasal_Cartilage|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C300|Nasal_Cartilage|882|Sarcoma|8825/3|Sarcoma
C300|Nasal_Cartilage|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C300|Nasal_Cartilage|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C300|Nasal_Cartilage|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C300|Nasal_Cartilage|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C300|Nasal_Cartilage|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C300|Nasal_Cartilage|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C300|Nasal_Cartilage|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C300|Nasal_Cartilage|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C300|Nasal_Cartilage|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C300|Nasal_Cartilage|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C300|Nasal_Cartilage|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C300|Nasal_Cartilage|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C300|Nasal_Cartilage|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C300|Nasal_Cartilage|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C300|Nasal_Cartilage|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C300|Nasal_Cartilage|904|Synovial_Sarcoma|9045/3|Sarcoma
C300|Nasal_Cartilage|922|Chondrosarcoma|9220/3|Chondrosarcoma
C300|Nasal_Cartilage|922|Chondrosarcoma|9221/3|Periosteal_Chondrosarcoma
C300|Nasal_Cartilage|937|Chordoma|9370/3|Chordoma
C300|Nasal_Cartilage|937|Chordoma|9371/3|Chondroid_Chordoma
C300|Nasal_Cartilage|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C300|Nasal_Cartilage|950|Neuroblastoma|9500/3|Neuroblastoma
C300|Nasal_Cartilage|950|Neuroblastoma|9501/3|Medulloepithelioma
C300|Nasal_Cartilage|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C300|Nasal_Cartilage|950|Neuroblastoma|9503/3|Neuroepithelioma
C300|Nasal_Cartilage|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C300|Nasal_Cartilage|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C300|Nasal_Cartilage|952|Neoplasm|9520/3|Neoplasm
C300|Nasal_Cartilage|952|Neoplasm|9521/3|Olfactory_Neurocytoma
C300|Nasal_Cartilage|952|Neoplasm|9522/3|Olfactory_Neuroblastoma
C300|Nasal_Cartilage|952|Neoplasm|9523/3|Olfactory_Neuroblastoma
C300|Nasal_Cartilage|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C300|Nasal_Cartilage|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C300|Nasal_Cartilage|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C300|Nasal_Cartilage|959|Lymphoma|9590/3|Lymphoma
C300|Nasal_Cartilage|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C300|Nasal_Cartilage|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C300|Nasal_Cartilage|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C300|Nasal_Cartilage|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C300|Nasal_Cartilage|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C300|Nasal_Cartilage|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C300|Nasal_Cartilage|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C300|Nasal_Cartilage|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C300|Nasal_Cartilage|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C300|Nasal_Cartilage|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C300|Nasal_Cartilage|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C300|Nasal_Cartilage|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C300|Nasal_Cartilage|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C300|Nasal_Cartilage|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C300|Nasal_Cartilage|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C300|Nasal_Cartilage|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C300|Nasal_Cartilage|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C300|Nasal_Cartilage|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C300|Nasal_Cartilage|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C300|Nasal_Cartilage|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C300|Nasal_Cartilage|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C300|Nasal_Cartilage|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C300|Nasal_Cartilage|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C300|Nasal_Cartilage|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C300|Nasal_Cartilage|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C300|Nasal_Cartilage|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C300|Nasal_Cartilage|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C300|Nasal_Cartilage|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C300|Nasal_Cartilage|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C300|Nasal_Cartilage|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C300|Nasal_Cartilage|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C300|Nasal_Cartilage|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C300|Nasal_Cartilage|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C300|Nasal_Cartilage|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C300|Nasal_Cartilage|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C300|Nasal_Cartilage|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C300|Nasal_Cartilage|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C300|Nasal_Cartilage|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C300|Nasal_Cartilage|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C300|Nasal_Cartilage|973|Plasmacytoma|9731/3|Plasmacytoma
C300|Nasal_Cartilage|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C300|Nasal_Cartilage|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C300|Nasal_Cartilage|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C300|Nasal_Cartilage|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C300|Nasal_Cartilage|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C300|Nasal_Cartilage|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C300|Nasal_Cartilage|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C300|Nasal_Cartilage|975|Neoplasm|9750/3|Malignant_Histiocytosis
C300|Nasal_Cartilage|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C300|Nasal_Cartilage|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C300|Nasal_Cartilage|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C300|Nasal_Cartilage|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C300|Nasal_Cartilage|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C300|Nasal_Cartilage|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C300|Nasal_Cartilage|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C300|Nasal_Cartilage|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C300|Nasal_Cartilage|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C300|Nasal_Cartilage|981|Neoplasm|9812/3|Lymphoma
C300|Nasal_Cartilage|981|Neoplasm|9813/3|Lymphoma
C300|Nasal_Cartilage|981|Neoplasm|9814/3|Lymphoma
C300|Nasal_Cartilage|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C300|Nasal_Cartilage|981|Neoplasm|9816/3|Hypodiploid_ALL
C300|Nasal_Cartilage|981|Neoplasm|9817/3|Lymphoma
C300|Nasal_Cartilage|981|Neoplasm|9818/3|Lymphoma
C300|Nasal_Cartilage|981|Neoplasm|9819/3|Leukemia__B_Cell
C300|Nasal_Cartilage|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C300|Nasal_Cartilage|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C300|Nasal_Cartilage|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C300|Nasal_Cartilage|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C300|Nasal_Cartilage|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C300|Nasal_Cartilage|997|Neoplasm|9971/3|Polymorphic_PTLD
C300|Nasal_Cartilage|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C301|Middle_Ear|800|Neoplasm|8000/3|Malignant_Neoplasm
C301|Middle_Ear|800|Neoplasm|8001/3|Malignant_Cell
C301|Middle_Ear|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C301|Middle_Ear|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C301|Middle_Ear|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C301|Middle_Ear|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C301|Middle_Ear|801|Carcinoma|8010/2|In_Situ_Cancer
C301|Middle_Ear|801|Carcinoma|8010/3|Carcinoma
C301|Middle_Ear|801|Carcinoma|8011/3|Malignant_Epithelioma
C301|Middle_Ear|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C301|Middle_Ear|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C301|Middle_Ear|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C301|Middle_Ear|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C301|Middle_Ear|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C301|Middle_Ear|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C301|Middle_Ear|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C301|Middle_Ear|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C301|Middle_Ear|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C301|Middle_Ear|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C301|Middle_Ear|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C301|Middle_Ear|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C301|Middle_Ear|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C301|Middle_Ear|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C301|Middle_Ear|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C301|Middle_Ear|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C301|Middle_Ear|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C301|Middle_Ear|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C301|Middle_Ear|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C301|Middle_Ear|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C301|Middle_Ear|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C301|Middle_Ear|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C301|Middle_Ear|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C301|Middle_Ear|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C301|Middle_Ear|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C301|Middle_Ear|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C301|Middle_Ear|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C301|Middle_Ear|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C301|Middle_Ear|813|Carcinoma|8130/2|Carcinoma
C301|Middle_Ear|813|Carcinoma|8130/3|Carcinoma
C301|Middle_Ear|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C301|Middle_Ear|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C301|Middle_Ear|814|Adenocarcinoma|8140/3|Adenocarcinoma
C301|Middle_Ear|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C301|Middle_Ear|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C301|Middle_Ear|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C301|Middle_Ear|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C301|Middle_Ear|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C301|Middle_Ear|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C301|Middle_Ear|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C301|Middle_Ear|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C301|Middle_Ear|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C301|Middle_Ear|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C301|Middle_Ear|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C301|Middle_Ear|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C301|Middle_Ear|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C301|Middle_Ear|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C301|Middle_Ear|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C301|Middle_Ear|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C301|Middle_Ear|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C301|Middle_Ear|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C301|Middle_Ear|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C301|Middle_Ear|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C301|Middle_Ear|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C301|Middle_Ear|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C301|Middle_Ear|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C301|Middle_Ear|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C301|Middle_Ear|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C301|Middle_Ear|872|Melanoma|8720/3|Melanoma
C301|Middle_Ear|872|Melanoma|8721/3|Nodular_Melanoma
C301|Middle_Ear|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C301|Middle_Ear|872|Melanoma|8723/3|Regressing_Melanoma
C301|Middle_Ear|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C301|Middle_Ear|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C301|Middle_Ear|874|Nevus|8745/3|Desmoplastic_Melanoma
C301|Middle_Ear|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C301|Middle_Ear|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C301|Middle_Ear|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C301|Middle_Ear|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C301|Middle_Ear|880|Sarcoma|8800/3|Sarcoma
C301|Middle_Ear|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C301|Middle_Ear|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C301|Middle_Ear|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C301|Middle_Ear|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C301|Middle_Ear|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C301|Middle_Ear|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C301|Middle_Ear|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C301|Middle_Ear|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C301|Middle_Ear|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C301|Middle_Ear|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C301|Middle_Ear|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C301|Middle_Ear|882|Sarcoma|8825/3|Sarcoma
C301|Middle_Ear|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C301|Middle_Ear|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C301|Middle_Ear|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C301|Middle_Ear|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C301|Middle_Ear|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C301|Middle_Ear|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C301|Middle_Ear|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C301|Middle_Ear|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C301|Middle_Ear|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C301|Middle_Ear|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C301|Middle_Ear|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C301|Middle_Ear|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C301|Middle_Ear|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C301|Middle_Ear|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C301|Middle_Ear|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C301|Middle_Ear|937|Chordoma|9370/3|Chordoma
C301|Middle_Ear|937|Chordoma|9371/3|Chondroid_Chordoma
C301|Middle_Ear|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C301|Middle_Ear|950|Neuroblastoma|9500/3|Neuroblastoma
C301|Middle_Ear|950|Neuroblastoma|9501/3|Medulloepithelioma
C301|Middle_Ear|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C301|Middle_Ear|950|Neuroblastoma|9503/3|Neuroepithelioma
C301|Middle_Ear|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C301|Middle_Ear|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C301|Middle_Ear|952|Neoplasm|9520/3|Neoplasm
C301|Middle_Ear|952|Neoplasm|9521/3|Olfactory_Neurocytoma
C301|Middle_Ear|952|Neoplasm|9522/3|Olfactory_Neuroblastoma
C301|Middle_Ear|952|Neoplasm|9523/3|Olfactory_Neuroblastoma
C301|Middle_Ear|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C301|Middle_Ear|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C301|Middle_Ear|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C301|Middle_Ear|957|Perineurioma|9571/3|Malignant_Perineurioma
C301|Middle_Ear|959|Lymphoma|9590/3|Lymphoma
C301|Middle_Ear|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C301|Middle_Ear|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C301|Middle_Ear|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C301|Middle_Ear|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C301|Middle_Ear|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C301|Middle_Ear|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C301|Middle_Ear|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C301|Middle_Ear|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C301|Middle_Ear|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C301|Middle_Ear|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C301|Middle_Ear|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C301|Middle_Ear|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C301|Middle_Ear|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C301|Middle_Ear|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C301|Middle_Ear|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C301|Middle_Ear|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C301|Middle_Ear|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C301|Middle_Ear|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C301|Middle_Ear|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C301|Middle_Ear|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C301|Middle_Ear|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C301|Middle_Ear|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C301|Middle_Ear|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C301|Middle_Ear|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C301|Middle_Ear|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C301|Middle_Ear|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C301|Middle_Ear|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C301|Middle_Ear|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C301|Middle_Ear|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C301|Middle_Ear|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C301|Middle_Ear|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C301|Middle_Ear|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C301|Middle_Ear|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C301|Middle_Ear|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C301|Middle_Ear|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C301|Middle_Ear|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C301|Middle_Ear|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C301|Middle_Ear|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C301|Middle_Ear|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C301|Middle_Ear|973|Plasmacytoma|9731/3|Plasmacytoma
C301|Middle_Ear|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C301|Middle_Ear|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C301|Middle_Ear|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C301|Middle_Ear|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C301|Middle_Ear|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C301|Middle_Ear|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C301|Middle_Ear|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C301|Middle_Ear|975|Neoplasm|9750/3|Malignant_Histiocytosis
C301|Middle_Ear|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C301|Middle_Ear|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C301|Middle_Ear|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C301|Middle_Ear|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C301|Middle_Ear|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C301|Middle_Ear|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C301|Middle_Ear|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C301|Middle_Ear|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C301|Middle_Ear|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C301|Middle_Ear|981|Neoplasm|9812/3|Lymphoma
C301|Middle_Ear|981|Neoplasm|9813/3|Lymphoma
C301|Middle_Ear|981|Neoplasm|9814/3|Lymphoma
C301|Middle_Ear|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C301|Middle_Ear|981|Neoplasm|9816/3|Hypodiploid_ALL
C301|Middle_Ear|981|Neoplasm|9817/3|Lymphoma
C301|Middle_Ear|981|Neoplasm|9818/3|Lymphoma
C301|Middle_Ear|981|Neoplasm|9819/3|Leukemia__B_Cell
C301|Middle_Ear|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C301|Middle_Ear|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C301|Middle_Ear|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C301|Middle_Ear|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C301|Middle_Ear|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C301|Middle_Ear|997|Neoplasm|9971/3|Polymorphic_PTLD
C301|Middle_Ear|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C310-C313, C318|Nasal_Sinus|800|Neoplasm|8000/3|Malignant_Neoplasm
C310-C313, C318|Nasal_Sinus|800|Neoplasm|8001/3|Malignant_Cell
C310-C313, C318|Nasal_Sinus|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C310-C313, C318|Nasal_Sinus|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C310-C313, C318|Nasal_Sinus|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C310-C313, C318|Nasal_Sinus|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C310-C313, C318|Nasal_Sinus|801|Carcinoma|8010/2|In_Situ_Cancer
C310-C313, C318|Nasal_Sinus|801|Carcinoma|8010/3|Carcinoma
C310-C313, C318|Nasal_Sinus|801|Carcinoma|8011/3|Malignant_Epithelioma
C310-C313, C318|Nasal_Sinus|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C310-C313, C318|Nasal_Sinus|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C310-C313, C318|Nasal_Sinus|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C310-C313, C318|Nasal_Sinus|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C310-C313, C318|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C310-C313, C318|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C310-C313, C318|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C310-C313, C318|Nasal_Sinus|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C310-C313, C318|Nasal_Sinus|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C310-C313, C318|Nasal_Sinus|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C310-C313, C318|Nasal_Sinus|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C310-C313, C318|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C310-C313, C318|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8085/3|Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8086/3|Squamous_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C310-C313, C318|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C310-C313, C318|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C310-C313, C318|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C310-C313, C318|Nasal_Sinus|813|Carcinoma|8130/2|Carcinoma
C310-C313, C318|Nasal_Sinus|813|Carcinoma|8130/3|Carcinoma
C310-C313, C318|Nasal_Sinus|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C310-C313, C318|Nasal_Sinus|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C310-C313, C318|Nasal_Sinus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C310-C313, C318|Nasal_Sinus|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C310-C313, C318|Nasal_Sinus|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C310-C313, C318|Nasal_Sinus|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C310-C313, C318|Nasal_Sinus|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C310-C313, C318|Nasal_Sinus|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C310-C313, C318|Nasal_Sinus|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C310-C313, C318|Nasal_Sinus|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C310-C313, C318|Nasal_Sinus|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C310-C313, C318|Nasal_Sinus|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C310-C313, C318|Nasal_Sinus|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C310-C313, C318|Nasal_Sinus|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C310-C313, C318|Nasal_Sinus|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C310-C313, C318|Nasal_Sinus|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C310-C313, C318|Nasal_Sinus|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C310-C313, C318|Nasal_Sinus|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C310-C313, C318|Nasal_Sinus|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C310-C313, C318|Nasal_Sinus|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C310-C313, C318|Nasal_Sinus|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C310-C313, C318|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C310-C313, C318|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C310-C313, C318|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C310-C313, C318|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C310-C313, C318|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C310-C313, C318|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C310-C313, C318|Nasal_Sinus|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C310-C313, C318|Nasal_Sinus|872|Melanoma|8720/3|Melanoma
C310-C313, C318|Nasal_Sinus|872|Melanoma|8721/3|Nodular_Melanoma
C310-C313, C318|Nasal_Sinus|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C310-C313, C318|Nasal_Sinus|872|Melanoma|8723/3|Regressing_Melanoma
C310-C313, C318|Nasal_Sinus|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C310-C313, C318|Nasal_Sinus|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C310-C313, C318|Nasal_Sinus|874|Nevus|8745/3|Desmoplastic_Melanoma
C310-C313, C318|Nasal_Sinus|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C310-C313, C318|Nasal_Sinus|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C310-C313, C318|Nasal_Sinus|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C310-C313, C318|Nasal_Sinus|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C310-C313, C318|Nasal_Sinus|880|Sarcoma|8800/3|Sarcoma
C310-C313, C318|Nasal_Sinus|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C310-C313, C318|Nasal_Sinus|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C310-C313, C318|Nasal_Sinus|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C310-C313, C318|Nasal_Sinus|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C310-C313, C318|Nasal_Sinus|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C310-C313, C318|Nasal_Sinus|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C310-C313, C318|Nasal_Sinus|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C310-C313, C318|Nasal_Sinus|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C310-C313, C318|Nasal_Sinus|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C310-C313, C318|Nasal_Sinus|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C310-C313, C318|Nasal_Sinus|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C310-C313, C318|Nasal_Sinus|882|Sarcoma|8825/3|Sarcoma
C310-C313, C318|Nasal_Sinus|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C310-C313, C318|Nasal_Sinus|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C310-C313, C318|Nasal_Sinus|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C310-C313, C318|Nasal_Sinus|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C310-C313, C318|Nasal_Sinus|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C310-C313, C318|Nasal_Sinus|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C310-C313, C318|Nasal_Sinus|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C310-C313, C318|Nasal_Sinus|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C310-C313, C318|Nasal_Sinus|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C310-C313, C318|Nasal_Sinus|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C310-C313, C318|Nasal_Sinus|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C310-C313, C318|Nasal_Sinus|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C310-C313, C318|Nasal_Sinus|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C310-C313, C318|Nasal_Sinus|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C310-C313, C318|Nasal_Sinus|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C310-C313, C318|Nasal_Sinus|904|Synovial_Sarcoma|9045/3|Sarcoma
C310-C313, C318|Nasal_Sinus|937|Chordoma|9370/3|Chordoma
C310-C313, C318|Nasal_Sinus|937|Chordoma|9371/3|Chondroid_Chordoma
C310-C313, C318|Nasal_Sinus|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C310-C313, C318|Nasal_Sinus|950|Neuroblastoma|9500/3|Neuroblastoma
C310-C313, C318|Nasal_Sinus|950|Neuroblastoma|9501/3|Medulloepithelioma
C310-C313, C318|Nasal_Sinus|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C310-C313, C318|Nasal_Sinus|950|Neuroblastoma|9503/3|Neuroepithelioma
C310-C313, C318|Nasal_Sinus|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C310-C313, C318|Nasal_Sinus|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C310-C313, C318|Nasal_Sinus|952|Neoplasm|9520/3|Neoplasm
C310-C313, C318|Nasal_Sinus|952|Neoplasm|9521/3|Olfactory_Neurocytoma
C310-C313, C318|Nasal_Sinus|952|Neoplasm|9522/3|Olfactory_Neuroblastoma
C310-C313, C318|Nasal_Sinus|952|Neoplasm|9523/3|Olfactory_Neuroblastoma
C310-C313, C318|Nasal_Sinus|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C310-C313, C318|Nasal_Sinus|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C310-C313, C318|Nasal_Sinus|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C310-C313, C318|Nasal_Sinus|957|Perineurioma|9571/3|Malignant_Perineurioma
C310-C313, C318|Nasal_Sinus|959|Lymphoma|9590/3|Lymphoma
C310-C313, C318|Nasal_Sinus|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C310-C313, C318|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C310-C313, C318|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C310-C313, C318|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C310-C313, C318|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C310-C313, C318|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C310-C313, C318|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C310-C313, C318|Nasal_Sinus|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C310-C313, C318|Nasal_Sinus|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C310-C313, C318|Nasal_Sinus|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C310-C313, C318|Nasal_Sinus|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C310-C313, C318|Nasal_Sinus|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C310-C313, C318|Nasal_Sinus|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C310-C313, C318|Nasal_Sinus|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C310-C313, C318|Nasal_Sinus|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C310-C313, C318|Nasal_Sinus|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C310-C313, C318|Nasal_Sinus|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C310-C313, C318|Nasal_Sinus|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C310-C313, C318|Nasal_Sinus|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C310-C313, C318|Nasal_Sinus|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C310-C313, C318|Nasal_Sinus|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C310-C313, C318|Nasal_Sinus|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C310-C313, C318|Nasal_Sinus|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C310-C313, C318|Nasal_Sinus|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C310-C313, C318|Nasal_Sinus|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C310-C313, C318|Nasal_Sinus|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C310-C313, C318|Nasal_Sinus|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C310-C313, C318|Nasal_Sinus|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C310-C313, C318|Nasal_Sinus|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C310-C313, C318|Nasal_Sinus|973|Plasmacytoma|9731/3|Plasmacytoma
C310-C313, C318|Nasal_Sinus|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C310-C313, C318|Nasal_Sinus|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C310-C313, C318|Nasal_Sinus|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C310-C313, C318|Nasal_Sinus|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C310-C313, C318|Nasal_Sinus|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C310-C313, C318|Nasal_Sinus|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C310-C313, C318|Nasal_Sinus|975|Neoplasm|9750/3|Malignant_Histiocytosis
C310-C313, C318|Nasal_Sinus|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C310-C313, C318|Nasal_Sinus|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C310-C313, C318|Nasal_Sinus|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C310-C313, C318|Nasal_Sinus|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C310-C313, C318|Nasal_Sinus|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C310-C313, C318|Nasal_Sinus|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C310-C313, C318|Nasal_Sinus|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C310-C313, C318|Nasal_Sinus|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9812/3|Lymphoma
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9813/3|Lymphoma
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9814/3|Lymphoma
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9816/3|Hypodiploid_ALL
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9817/3|Lymphoma
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9818/3|Lymphoma
C310-C313, C318|Nasal_Sinus|981|Neoplasm|9819/3|Leukemia__B_Cell
C310-C313, C318|Nasal_Sinus|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C310-C313, C318|Nasal_Sinus|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C310-C313, C318|Nasal_Sinus|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C310-C313, C318|Nasal_Sinus|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C310-C313, C318|Nasal_Sinus|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C310-C313, C318|Nasal_Sinus|997|Neoplasm|9971/3|Polymorphic_PTLD
C310-C313, C318|Nasal_Sinus|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C319|Nasal_Sinus|800|Neoplasm|8000/3|Malignant_Neoplasm
C319|Nasal_Sinus|800|Neoplasm|8001/3|Malignant_Cell
C319|Nasal_Sinus|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C319|Nasal_Sinus|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C319|Nasal_Sinus|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C319|Nasal_Sinus|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C319|Nasal_Sinus|801|Carcinoma|8010/2|In_Situ_Cancer
C319|Nasal_Sinus|801|Carcinoma|8010/3|Carcinoma
C319|Nasal_Sinus|801|Carcinoma|8011/3|Malignant_Epithelioma
C319|Nasal_Sinus|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C319|Nasal_Sinus|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C319|Nasal_Sinus|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C319|Nasal_Sinus|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C319|Nasal_Sinus|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C319|Nasal_Sinus|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C319|Nasal_Sinus|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C319|Nasal_Sinus|802|Carcinoma|8023/3|NUT_Carcinoma
C319|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C319|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C319|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C319|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C319|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C319|Nasal_Sinus|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C319|Nasal_Sinus|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C319|Nasal_Sinus|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C319|Nasal_Sinus|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C319|Nasal_Sinus|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C319|Nasal_Sinus|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C319|Nasal_Sinus|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C319|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C319|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C319|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C319|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8085/3|Squamous_Cell_Carcinoma
C319|Nasal_Sinus|808|Lymphoepithelial_Carcinoma|8086/3|Squamous_Cell_Carcinoma
C319|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C319|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C319|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C319|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C319|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C319|Nasal_Sinus|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C319|Nasal_Sinus|813|Carcinoma|8130/2|Carcinoma
C319|Nasal_Sinus|813|Carcinoma|8130/3|Carcinoma
C319|Nasal_Sinus|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C319|Nasal_Sinus|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C319|Nasal_Sinus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C319|Nasal_Sinus|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C319|Nasal_Sinus|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C319|Nasal_Sinus|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C319|Nasal_Sinus|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C319|Nasal_Sinus|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C319|Nasal_Sinus|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C319|Nasal_Sinus|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C319|Nasal_Sinus|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C319|Nasal_Sinus|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C319|Nasal_Sinus|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C319|Nasal_Sinus|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C319|Nasal_Sinus|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C319|Nasal_Sinus|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C319|Nasal_Sinus|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C319|Nasal_Sinus|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C319|Nasal_Sinus|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C319|Nasal_Sinus|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C319|Nasal_Sinus|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C319|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C319|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C319|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C319|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C319|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C319|Nasal_Sinus|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C319|Nasal_Sinus|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C319|Nasal_Sinus|872|Melanoma|8720/3|Melanoma
C319|Nasal_Sinus|872|Melanoma|8721/3|Nodular_Melanoma
C319|Nasal_Sinus|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C319|Nasal_Sinus|872|Melanoma|8723/3|Regressing_Melanoma
C319|Nasal_Sinus|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C319|Nasal_Sinus|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C319|Nasal_Sinus|874|Nevus|8745/3|Desmoplastic_Melanoma
C319|Nasal_Sinus|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C319|Nasal_Sinus|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C319|Nasal_Sinus|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C319|Nasal_Sinus|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C319|Nasal_Sinus|880|Sarcoma|8800/3|Sarcoma
C319|Nasal_Sinus|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C319|Nasal_Sinus|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C319|Nasal_Sinus|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C319|Nasal_Sinus|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C319|Nasal_Sinus|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C319|Nasal_Sinus|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C319|Nasal_Sinus|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C319|Nasal_Sinus|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C319|Nasal_Sinus|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C319|Nasal_Sinus|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C319|Nasal_Sinus|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C319|Nasal_Sinus|882|Sarcoma|8825/3|Sarcoma
C319|Nasal_Sinus|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C319|Nasal_Sinus|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C319|Nasal_Sinus|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C319|Nasal_Sinus|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C319|Nasal_Sinus|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C319|Nasal_Sinus|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C319|Nasal_Sinus|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C319|Nasal_Sinus|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C319|Nasal_Sinus|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C319|Nasal_Sinus|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C319|Nasal_Sinus|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C319|Nasal_Sinus|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C319|Nasal_Sinus|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C319|Nasal_Sinus|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C319|Nasal_Sinus|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C319|Nasal_Sinus|904|Synovial_Sarcoma|9045/3|Sarcoma
C319|Nasal_Sinus|937|Chordoma|9370/3|Chordoma
C319|Nasal_Sinus|937|Chordoma|9371/3|Chondroid_Chordoma
C319|Nasal_Sinus|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C319|Nasal_Sinus|950|Neuroblastoma|9500/3|Neuroblastoma
C319|Nasal_Sinus|950|Neuroblastoma|9501/3|Medulloepithelioma
C319|Nasal_Sinus|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C319|Nasal_Sinus|950|Neuroblastoma|9503/3|Neuroepithelioma
C319|Nasal_Sinus|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C319|Nasal_Sinus|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C319|Nasal_Sinus|952|Neoplasm|9520/3|Neoplasm
C319|Nasal_Sinus|952|Neoplasm|9521/3|Olfactory_Neurocytoma
C319|Nasal_Sinus|952|Neoplasm|9522/3|Olfactory_Neuroblastoma
C319|Nasal_Sinus|952|Neoplasm|9523/3|Olfactory_Neuroblastoma
C319|Nasal_Sinus|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C319|Nasal_Sinus|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C319|Nasal_Sinus|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C319|Nasal_Sinus|957|Perineurioma|9571/3|Malignant_Perineurioma
C319|Nasal_Sinus|959|Lymphoma|9590/3|Lymphoma
C319|Nasal_Sinus|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C319|Nasal_Sinus|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C319|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C319|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C319|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C319|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C319|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C319|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C319|Nasal_Sinus|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C319|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C319|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C319|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C319|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C319|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C319|Nasal_Sinus|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C319|Nasal_Sinus|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C319|Nasal_Sinus|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C319|Nasal_Sinus|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C319|Nasal_Sinus|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C319|Nasal_Sinus|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C319|Nasal_Sinus|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C319|Nasal_Sinus|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C319|Nasal_Sinus|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C319|Nasal_Sinus|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C319|Nasal_Sinus|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C319|Nasal_Sinus|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C319|Nasal_Sinus|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C319|Nasal_Sinus|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C319|Nasal_Sinus|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C319|Nasal_Sinus|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C319|Nasal_Sinus|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C319|Nasal_Sinus|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C319|Nasal_Sinus|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C319|Nasal_Sinus|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C319|Nasal_Sinus|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C319|Nasal_Sinus|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C319|Nasal_Sinus|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C319|Nasal_Sinus|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C319|Nasal_Sinus|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C319|Nasal_Sinus|973|Plasmacytoma|9731/3|Plasmacytoma
C319|Nasal_Sinus|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C319|Nasal_Sinus|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C319|Nasal_Sinus|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C319|Nasal_Sinus|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C319|Nasal_Sinus|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C319|Nasal_Sinus|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C319|Nasal_Sinus|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C319|Nasal_Sinus|975|Neoplasm|9750/3|Malignant_Histiocytosis
C319|Nasal_Sinus|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C319|Nasal_Sinus|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C319|Nasal_Sinus|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C319|Nasal_Sinus|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C319|Nasal_Sinus|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C319|Nasal_Sinus|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C319|Nasal_Sinus|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C319|Nasal_Sinus|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C319|Nasal_Sinus|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C319|Nasal_Sinus|981|Neoplasm|9812/3|Lymphoma
C319|Nasal_Sinus|981|Neoplasm|9813/3|Lymphoma
C319|Nasal_Sinus|981|Neoplasm|9814/3|Lymphoma
C319|Nasal_Sinus|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C319|Nasal_Sinus|981|Neoplasm|9816/3|Hypodiploid_ALL
C319|Nasal_Sinus|981|Neoplasm|9817/3|Lymphoma
C319|Nasal_Sinus|981|Neoplasm|9818/3|Lymphoma
C319|Nasal_Sinus|981|Neoplasm|9819/3|Leukemia__B_Cell
C319|Nasal_Sinus|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C319|Nasal_Sinus|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C319|Nasal_Sinus|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C319|Nasal_Sinus|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C319|Nasal_Sinus|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C319|Nasal_Sinus|997|Neoplasm|9971/3|Polymorphic_PTLD
C319|Nasal_Sinus|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C320-C323,C328-C329|Larynx|800|Neoplasm|8000/3|Malignant_Neoplasm
C320-C323,C328-C329|Larynx|800|Neoplasm|8001/3|Malignant_Cell
C320-C323,C328-C329|Larynx|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C320-C323,C328-C329|Larynx|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C320-C323,C328-C329|Larynx|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C320-C323,C328-C329|Larynx|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C320-C323,C328-C329|Larynx|801|Carcinoma|8010/2|In_Situ_Cancer
C320-C323,C328-C329|Larynx|801|Carcinoma|8010/3|Carcinoma
C320-C323,C328-C329|Larynx|801|Carcinoma|8011/3|Malignant_Epithelioma
C320-C323,C328-C329|Larynx|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C320-C323,C328-C329|Larynx|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C320-C323,C328-C329|Larynx|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C320-C323,C328-C329|Larynx|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C320-C323,C328-C329|Larynx|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C320-C323,C328-C329|Larynx|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C320-C323,C328-C329|Larynx|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C320-C323,C328-C329|Larynx|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C320-C323,C328-C329|Larynx|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C320-C323,C328-C329|Larynx|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C320-C323,C328-C329|Larynx|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C320-C323,C328-C329|Larynx|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C320-C323,C328-C329|Larynx|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C320-C323,C328-C329|Larynx|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C320-C323,C328-C329|Larynx|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C320-C323,C328-C329|Larynx|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C320-C323,C328-C329|Larynx|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C320-C323,C328-C329|Larynx|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C320-C323,C328-C329|Larynx|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C320-C323,C328-C329|Larynx|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C320-C323,C328-C329|Larynx|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C320-C323,C328-C329|Larynx|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C320-C323,C328-C329|Larynx|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C320-C323,C328-C329|Larynx|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C320-C323,C328-C329|Larynx|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C320-C323,C328-C329|Larynx|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C320-C323,C328-C329|Larynx|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8140/3|Adenocarcinoma
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C320-C323,C328-C329|Larynx|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C320-C323,C328-C329|Larynx|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C320-C323,C328-C329|Larynx|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C320-C323,C328-C329|Larynx|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C320-C323,C328-C329|Larynx|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C320-C323,C328-C329|Larynx|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C320-C323,C328-C329|Larynx|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C320-C323,C328-C329|Larynx|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C320-C323,C328-C329|Larynx|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C320-C323,C328-C329|Larynx|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C320-C323,C328-C329|Larynx|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C320-C323,C328-C329|Larynx|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C320-C323,C328-C329|Larynx|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C320-C323,C328-C329|Larynx|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C320-C323,C328-C329|Larynx|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C320-C323,C328-C329|Larynx|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8800/3|Sarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C320-C323,C328-C329|Larynx|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C320-C323,C328-C329|Larynx|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C320-C323,C328-C329|Larynx|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C320-C323,C328-C329|Larynx|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C320-C323,C328-C329|Larynx|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C320-C323,C328-C329|Larynx|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C320-C323,C328-C329|Larynx|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C320-C323,C328-C329|Larynx|882|Sarcoma|8825/3|Sarcoma
C320-C323,C328-C329|Larynx|898|Carcinosarcoma|8980/3|Carcinosarcoma
C320-C323,C328-C329|Larynx|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C320-C323,C328-C329|Larynx|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C320-C323,C328-C329|Larynx|922|Chondrosarcoma|9220/3|Chondrosarcoma
C320-C323,C328-C329|Larynx|922|Chondrosarcoma|9221/3|Periosteal_Chondrosarcoma
C320-C323,C328-C329|Larynx|959|Lymphoma|9590/3|Lymphoma
C320-C323,C328-C329|Larynx|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C320-C323,C328-C329|Larynx|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C320-C323,C328-C329|Larynx|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C320-C323,C328-C329|Larynx|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C320-C323,C328-C329|Larynx|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C320-C323,C328-C329|Larynx|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C320-C323,C328-C329|Larynx|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C320-C323,C328-C329|Larynx|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C320-C323,C328-C329|Larynx|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C320-C323,C328-C329|Larynx|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C320-C323,C328-C329|Larynx|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C320-C323,C328-C329|Larynx|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C320-C323,C328-C329|Larynx|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C320-C323,C328-C329|Larynx|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C320-C323,C328-C329|Larynx|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C320-C323,C328-C329|Larynx|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C320-C323,C328-C329|Larynx|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C320-C323,C328-C329|Larynx|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C320-C323,C328-C329|Larynx|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C320-C323,C328-C329|Larynx|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C320-C323,C328-C329|Larynx|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C320-C323,C328-C329|Larynx|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C320-C323,C328-C329|Larynx|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C320-C323,C328-C329|Larynx|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C320-C323,C328-C329|Larynx|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C320-C323,C328-C329|Larynx|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C320-C323,C328-C329|Larynx|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C320-C323,C328-C329|Larynx|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C320-C323,C328-C329|Larynx|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9731/3|Plasmacytoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C320-C323,C328-C329|Larynx|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C320-C323,C328-C329|Larynx|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C320-C323,C328-C329|Larynx|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C320-C323,C328-C329|Larynx|975|Neoplasm|9750/3|Malignant_Histiocytosis
C320-C323,C328-C329|Larynx|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C320-C323,C328-C329|Larynx|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C320-C323,C328-C329|Larynx|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C320-C323,C328-C329|Larynx|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C320-C323,C328-C329|Larynx|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C320-C323,C328-C329|Larynx|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C320-C323,C328-C329|Larynx|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C320-C323,C328-C329|Larynx|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C320-C323,C328-C329|Larynx|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C320-C323,C328-C329|Larynx|981|Neoplasm|9812/3|Lymphoma
C320-C323,C328-C329|Larynx|981|Neoplasm|9813/3|Lymphoma
C320-C323,C328-C329|Larynx|981|Neoplasm|9814/3|Lymphoma
C320-C323,C328-C329|Larynx|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C320-C323,C328-C329|Larynx|981|Neoplasm|9816/3|Hypodiploid_ALL
C320-C323,C328-C329|Larynx|981|Neoplasm|9817/3|Lymphoma
C320-C323,C328-C329|Larynx|981|Neoplasm|9818/3|Lymphoma
C320-C323,C328-C329|Larynx|981|Neoplasm|9819/3|Leukemia__B_Cell
C320-C323,C328-C329|Larynx|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C320-C323,C328-C329|Larynx|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C320-C323,C328-C329|Larynx|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C320-C323,C328-C329|Larynx|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C320-C323,C328-C329|Larynx|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C320-C323,C328-C329|Larynx|997|Neoplasm|9971/3|Polymorphic_PTLD
C320-C323,C328-C329|Larynx|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C339|Trachea|800|Neoplasm|8000/3|Malignant_Neoplasm
C339|Trachea|800|Neoplasm|8001/3|Malignant_Cell
C339|Trachea|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C339|Trachea|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C339|Trachea|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C339|Trachea|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C339|Trachea|801|Carcinoma|8010/2|In_Situ_Cancer
C339|Trachea|801|Carcinoma|8010/3|Carcinoma
C339|Trachea|801|Carcinoma|8011/3|Malignant_Epithelioma
C339|Trachea|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C339|Trachea|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C339|Trachea|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C339|Trachea|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C339|Trachea|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C339|Trachea|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C339|Trachea|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C339|Trachea|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C339|Trachea|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C339|Trachea|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C339|Trachea|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C339|Trachea|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C339|Trachea|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C339|Trachea|804|Non_Small_Cell_Carcinoma|8046/3|Non_Small_Cell_Carcinoma
C339|Trachea|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C339|Trachea|804|Small_Cell_Carcinoma|8042/3|Small_Cell_Carcinoma
C339|Trachea|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C339|Trachea|804|Small_Cell_Carcinoma|8044/3|Small_Cell_Intermediate_Cell_Carcinoma
C339|Trachea|804|Small_Cell_Carcinoma|8045/3|Combined_Small_Cell_Lung_Carcinoma
C339|Trachea|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C339|Trachea|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C339|Trachea|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C339|Trachea|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C339|Trachea|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C339|Trachea|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C339|Trachea|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C339|Trachea|814|Adenocarcinoma|8140/3|Adenocarcinoma
C339|Trachea|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C339|Trachea|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C339|Trachea|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C339|Trachea|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C339|Trachea|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C339|Trachea|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C339|Trachea|825|Bronchioloalveolar_Adenocarcinoma|8250/3|null
C339|Trachea|825|Bronchioloalveolar_Adenocarcinoma|8252/3|Bronchioloalveolar_Adenocarcinoma
C339|Trachea|825|Bronchioloalveolar_Adenocarcinoma|8253/3|Mucinous_Adenocarcinoma
C339|Trachea|825|Bronchioloalveolar_Adenocarcinoma|8254/3|Adenocarcinoma
C339|Trachea|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C339|Trachea|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C339|Trachea|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C339|Trachea|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C339|Trachea|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C339|Trachea|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C339|Trachea|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C339|Trachea|880|Sarcoma|8800/3|Sarcoma
C339|Trachea|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C339|Trachea|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C339|Trachea|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C339|Trachea|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C339|Trachea|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C339|Trachea|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C339|Trachea|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C339|Trachea|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C339|Trachea|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C339|Trachea|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C339|Trachea|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C339|Trachea|882|Sarcoma|8825/3|Sarcoma
C339|Trachea|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C339|Trachea|897|Hepatoblastoma|8972/3|Pulmonary_Blastoma
C339|Trachea|897|Hepatoblastoma|8973/3|Pleuropulmonary_Blastoma
C339|Trachea|922|Chondrosarcoma|9220/3|Chondrosarcoma
C339|Trachea|922|Chondrosarcoma|9221/3|Periosteal_Chondrosarcoma
C339|Trachea|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C339|Trachea|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C340-C343,C348-C349|Bronchus|800|Neoplasm|8000/3|Malignant_Neoplasm
C340-C343,C348-C349|Bronchus|800|Neoplasm|8001/3|Malignant_Cell
C340-C343,C348-C349|Bronchus|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C340-C343,C348-C349|Bronchus|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C340-C343,C348-C349|Bronchus|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C340-C343,C348-C349|Bronchus|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C340-C343,C348-C349|Bronchus|801|Carcinoma|8010/2|In_Situ_Cancer
C340-C343,C348-C349|Bronchus|801|Carcinoma|8010/3|Carcinoma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8011/3|Malignant_Epithelioma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C340-C343,C348-C349|Bronchus|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C340-C343,C348-C349|Bronchus|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C340-C343,C348-C349|Bronchus|802|Carcinoma|8023/3|NUT_Carcinoma
C340-C343,C348-C349|Bronchus|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C340-C343,C348-C349|Bronchus|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C340-C343,C348-C349|Bronchus|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C340-C343,C348-C349|Bronchus|804|Non_Small_Cell_Carcinoma|8046/3|Non_Small_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|804|Small_Cell_Carcinoma|8042/3|Small_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C340-C343,C348-C349|Bronchus|804|Small_Cell_Carcinoma|8044/3|Small_Cell_Intermediate_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|804|Small_Cell_Carcinoma|8045/3|Combined_Small_Cell_Lung_Carcinoma
C340-C343,C348-C349|Bronchus|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C340-C343,C348-C349|Bronchus|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C340-C343,C348-C349|Bronchus|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C340-C343,C348-C349|Bronchus|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C340-C343,C348-C349|Bronchus|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C340-C343,C348-C349|Bronchus|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C340-C343,C348-C349|Bronchus|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C340-C343,C348-C349|Bronchus|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C340-C343,C348-C349|Bronchus|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C340-C343,C348-C349|Bronchus|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C340-C343,C348-C349|Bronchus|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C340-C343,C348-C349|Bronchus|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C340-C343,C348-C349|Bronchus|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C340-C343,C348-C349|Bronchus|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C340-C343,C348-C349|Bronchus|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C340-C343,C348-C349|Bronchus|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C340-C343,C348-C349|Bronchus|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C340-C343,C348-C349|Bronchus|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C340-C343,C348-C349|Bronchus|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C340-C343,C348-C349|Bronchus|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C340-C343,C348-C349|Bronchus|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C340-C343,C348-C349|Bronchus|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C340-C343,C348-C349|Bronchus|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8250/2|Adenocarcinoma_In_Situ
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8250/3|null
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8251/3|Bronchioloalveolar_Adenocarcinoma
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8252/3|Bronchioloalveolar_Adenocarcinoma
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8253/2|Adenocarcinoma_In_Situ
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8253/3|Mucinous_Adenocarcinoma
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8254/3|Adenocarcinoma
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8256/3|Adenocarcinoma
C340-C343,C348-C349|Bronchus|825|Bronchioloalveolar_Adenocarcinoma|8257/3|Mucinous_Adenocarcinoma
C340-C343,C348-C349|Bronchus|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C340-C343,C348-C349|Bronchus|826|Papillary_Adenocarcinoma|8265/3|Micropapillary_Carcinoma
C340-C343,C348-C349|Bronchus|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C340-C343,C348-C349|Bronchus|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C340-C343,C348-C349|Bronchus|833|Follicular_Thyroid_Carcinoma|8333/3|Fetal_Adenocarcinoma
C340-C343,C348-C349|Bronchus|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C340-C343,C348-C349|Bronchus|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C340-C343,C348-C349|Bronchus|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C340-C343,C348-C349|Bronchus|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C340-C343,C348-C349|Bronchus|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C340-C343,C348-C349|Bronchus|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C340-C343,C348-C349|Bronchus|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C340-C343,C348-C349|Bronchus|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C340-C343,C348-C349|Bronchus|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C340-C343,C348-C349|Bronchus|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C340-C343,C348-C349|Bronchus|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C340-C343,C348-C349|Bronchus|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C340-C343,C348-C349|Bronchus|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C340-C343,C348-C349|Bronchus|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C340-C343,C348-C349|Bronchus|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C340-C343,C348-C349|Bronchus|871|Malignant_Glomus_Tumor|8714/3|Malignant_PEComa
C340-C343,C348-C349|Bronchus|880|Sarcoma|8800/3|Sarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C340-C343,C348-C349|Bronchus|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C340-C343,C348-C349|Bronchus|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C340-C343,C348-C349|Bronchus|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C340-C343,C348-C349|Bronchus|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C340-C343,C348-C349|Bronchus|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C340-C343,C348-C349|Bronchus|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C340-C343,C348-C349|Bronchus|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C340-C343,C348-C349|Bronchus|882|Sarcoma|8825/3|Sarcoma
C340-C343,C348-C349|Bronchus|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C340-C343,C348-C349|Bronchus|884|Myxosarcoma|8842/3|Sarcoma
C340-C343,C348-C349|Bronchus|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C340-C343,C348-C349|Bronchus|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C340-C343,C348-C349|Bronchus|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C340-C343,C348-C349|Bronchus|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C340-C343,C348-C349|Bronchus|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C340-C343,C348-C349|Bronchus|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C340-C343,C348-C349|Bronchus|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C340-C343,C348-C349|Bronchus|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C340-C343,C348-C349|Bronchus|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C340-C343,C348-C349|Bronchus|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C340-C343,C348-C349|Bronchus|897|Hepatoblastoma|8972/3|Pulmonary_Blastoma
C340-C343,C348-C349|Bronchus|897|Hepatoblastoma|8973/3|Pleuropulmonary_Blastoma
C340-C343,C348-C349|Bronchus|898|Carcinosarcoma|8980/3|Carcinosarcoma
C340-C343,C348-C349|Bronchus|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C340-C343,C348-C349|Bronchus|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C340-C343,C348-C349|Bronchus|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C340-C343,C348-C349|Bronchus|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C340-C343,C348-C349|Bronchus|905|Malignant_Mesothelioma|9050/3|Malignant_Mesothelioma
C340-C343,C348-C349|Bronchus|905|Malignant_Mesothelioma|9051/3|Sarcomatoid_Mesothelioma
C340-C343,C348-C349|Bronchus|905|Malignant_Mesothelioma|9052/3|Mesothelioma
C340-C343,C348-C349|Bronchus|905|Malignant_Mesothelioma|9053/3|Biphasic_Mesothelioma
C340-C343,C348-C349|Bronchus|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C340-C343,C348-C349|Bronchus|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C340-C343,C348-C349|Bronchus|913|Hemangioendothelioma|9137/3|Intimal_Sarcoma
C340-C343,C348-C349|Bronchus|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C340-C343,C348-C349|Bronchus|959|Lymphoma|9590/3|Lymphoma
C340-C343,C348-C349|Bronchus|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C340-C343,C348-C349|Bronchus|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C340-C343,C348-C349|Bronchus|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C340-C343,C348-C349|Bronchus|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C340-C343,C348-C349|Bronchus|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C340-C343,C348-C349|Bronchus|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C340-C343,C348-C349|Bronchus|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C340-C343,C348-C349|Bronchus|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C340-C343,C348-C349|Bronchus|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C340-C343,C348-C349|Bronchus|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C340-C343,C348-C349|Bronchus|967|B_Cell_Lymphomas|9678/3|Primary_Effusion_Lymphoma
C340-C343,C348-C349|Bronchus|967|B_Cell_Lymphomas|9679/3|Mediastinal_Large_B_cell_Lymphoma
C340-C343,C348-C349|Bronchus|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C340-C343,C348-C349|Bronchus|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C340-C343,C348-C349|Bronchus|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C340-C343,C348-C349|Bronchus|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C340-C343,C348-C349|Bronchus|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C340-C343,C348-C349|Bronchus|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C340-C343,C348-C349|Bronchus|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C340-C343,C348-C349|Bronchus|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C340-C343,C348-C349|Bronchus|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C340-C343,C348-C349|Bronchus|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C340-C343,C348-C349|Bronchus|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C340-C343,C348-C349|Bronchus|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C340-C343,C348-C349|Bronchus|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C340-C343,C348-C349|Bronchus|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C340-C343,C348-C349|Bronchus|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C340-C343,C348-C349|Bronchus|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C340-C343,C348-C349|Bronchus|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C340-C343,C348-C349|Bronchus|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C340-C343,C348-C349|Bronchus|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9731/3|Plasmacytoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C340-C343,C348-C349|Bronchus|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C340-C343,C348-C349|Bronchus|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C340-C343,C348-C349|Bronchus|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C340-C343,C348-C349|Bronchus|975|Neoplasm|9750/3|Malignant_Histiocytosis
C340-C343,C348-C349|Bronchus|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C340-C343,C348-C349|Bronchus|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C340-C343,C348-C349|Bronchus|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C340-C343,C348-C349|Bronchus|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C340-C343,C348-C349|Bronchus|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C340-C343,C348-C349|Bronchus|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C340-C343,C348-C349|Bronchus|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C340-C343,C348-C349|Bronchus|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C340-C343,C348-C349|Bronchus|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C340-C343,C348-C349|Bronchus|981|Neoplasm|9812/3|Lymphoma
C340-C343,C348-C349|Bronchus|981|Neoplasm|9813/3|Lymphoma
C340-C343,C348-C349|Bronchus|981|Neoplasm|9814/3|Lymphoma
C340-C343,C348-C349|Bronchus|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C340-C343,C348-C349|Bronchus|981|Neoplasm|9816/3|Hypodiploid_ALL
C340-C343,C348-C349|Bronchus|981|Neoplasm|9817/3|Lymphoma
C340-C343,C348-C349|Bronchus|981|Neoplasm|9818/3|Lymphoma
C340-C343,C348-C349|Bronchus|981|Neoplasm|9819/3|Leukemia__B_Cell
C340-C343,C348-C349|Bronchus|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C340-C343,C348-C349|Bronchus|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C340-C343,C348-C349|Bronchus|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C340-C343,C348-C349|Bronchus|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C340-C343,C348-C349|Bronchus|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C340-C343,C348-C349|Bronchus|997|Neoplasm|9971/3|Polymorphic_PTLD
C340-C343,C348-C349|Bronchus|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C379|Thymus_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C379|Thymus_Gland|800|Neoplasm|8001/3|Malignant_Cell
C379|Thymus_Gland|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C379|Thymus_Gland|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C379|Thymus_Gland|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C379|Thymus_Gland|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C379|Thymus_Gland|801|Carcinoma|8010/2|In_Situ_Cancer
C379|Thymus_Gland|801|Carcinoma|8010/3|Carcinoma
C379|Thymus_Gland|801|Carcinoma|8011/3|Malignant_Epithelioma
C379|Thymus_Gland|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C379|Thymus_Gland|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C379|Thymus_Gland|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C379|Thymus_Gland|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C379|Thymus_Gland|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C379|Thymus_Gland|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C379|Thymus_Gland|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C379|Thymus_Gland|802|Carcinoma|8023/3|NUT_Carcinoma
C379|Thymus_Gland|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C379|Thymus_Gland|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C379|Thymus_Gland|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C379|Thymus_Gland|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C379|Thymus_Gland|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C379|Thymus_Gland|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C379|Thymus_Gland|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C379|Thymus_Gland|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C379|Thymus_Gland|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C379|Thymus_Gland|858|Malignant_Thymoma|8580/3|Malignant_Thymoma
C379|Thymus_Gland|858|Malignant_Thymoma|8581/3|Malignant_Type_A_Thymoma
C379|Thymus_Gland|858|Malignant_Thymoma|8582/3|Malignant_Type_AB_Thymoma
C379|Thymus_Gland|858|Malignant_Thymoma|8583/3|Malignant_Type_B1_Thymoma
C379|Thymus_Gland|858|Malignant_Thymoma|8584/3|Malignant_Type_B2_Thymoma
C379|Thymus_Gland|858|Malignant_Thymoma|8585/3|Thymoma_Type_B3
C379|Thymus_Gland|858|Malignant_Thymoma|8586/3|Thymic_Carcinoma
C379|Thymus_Gland|858|Malignant_Thymoma|8588/3|Neoplasm
C379|Thymus_Gland|858|Malignant_Thymoma|8589/3|Carcinoma_Showing_Thymus_like_Element
C379|Thymus_Gland|908|Teratoma|9086/3|Hematopoietic_Neoplasm
C379|Thymus_Gland|959|Lymphoma|9590/3|Lymphoma
C379|Thymus_Gland|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C379|Thymus_Gland|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C379|Thymus_Gland|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C379|Thymus_Gland|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C379|Thymus_Gland|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C379|Thymus_Gland|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C379|Thymus_Gland|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C379|Thymus_Gland|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C379|Thymus_Gland|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C379|Thymus_Gland|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C379|Thymus_Gland|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C379|Thymus_Gland|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C379|Thymus_Gland|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C379|Thymus_Gland|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C379|Thymus_Gland|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C379|Thymus_Gland|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C379|Thymus_Gland|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C379|Thymus_Gland|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C379|Thymus_Gland|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C379|Thymus_Gland|967|B_Cell_Lymphomas|9679/3|Mediastinal_Large_B_cell_Lymphoma
C379|Thymus_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C379|Thymus_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C379|Thymus_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C379|Thymus_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C379|Thymus_Gland|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C379|Thymus_Gland|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C379|Thymus_Gland|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C379|Thymus_Gland|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C379|Thymus_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C379|Thymus_Gland|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C379|Thymus_Gland|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C379|Thymus_Gland|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C379|Thymus_Gland|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C379|Thymus_Gland|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C379|Thymus_Gland|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C379|Thymus_Gland|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C379|Thymus_Gland|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C379|Thymus_Gland|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C379|Thymus_Gland|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C379|Thymus_Gland|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C379|Thymus_Gland|973|Plasmacytoma|9731/3|Plasmacytoma
C379|Thymus_Gland|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C379|Thymus_Gland|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C379|Thymus_Gland|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C379|Thymus_Gland|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C379|Thymus_Gland|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C379|Thymus_Gland|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C379|Thymus_Gland|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C379|Thymus_Gland|975|Neoplasm|9750/3|Malignant_Histiocytosis
C379|Thymus_Gland|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C379|Thymus_Gland|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C379|Thymus_Gland|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C379|Thymus_Gland|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C379|Thymus_Gland|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C379|Thymus_Gland|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C379|Thymus_Gland|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C379|Thymus_Gland|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C379|Thymus_Gland|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C379|Thymus_Gland|981|Neoplasm|9812/3|Lymphoma
C379|Thymus_Gland|981|Neoplasm|9813/3|Lymphoma
C379|Thymus_Gland|981|Neoplasm|9814/3|Lymphoma
C379|Thymus_Gland|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C379|Thymus_Gland|981|Neoplasm|9816/3|Hypodiploid_ALL
C379|Thymus_Gland|981|Neoplasm|9817/3|Lymphoma
C379|Thymus_Gland|981|Neoplasm|9818/3|Lymphoma
C379|Thymus_Gland|981|Neoplasm|9819/3|Leukemia__B_Cell
C379|Thymus_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C379|Thymus_Gland|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C379|Thymus_Gland|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C379|Thymus_Gland|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C379|Thymus_Gland|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C379|Thymus_Gland|997|Neoplasm|9971/3|Polymorphic_PTLD
C379|Thymus_Gland|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C380|Heart|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C380|Heart|913|Hemangioendothelioma|9137/3|Intimal_Sarcoma
C380|Heart|959|Lymphoma|9590/3|Lymphoma
C380|Heart|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C380|Heart|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C380|Heart|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C380|Heart|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C380|Heart|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C380|Heart|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C380|Heart|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C380|Heart|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C380|Heart|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C380|Heart|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C380|Heart|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C380|Heart|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C380|Heart|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C380|Heart|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C380|Heart|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C380|Heart|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C380|Heart|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C380|Heart|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C380|Heart|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C380|Heart|967|B_Cell_Lymphomas|9678/3|Primary_Effusion_Lymphoma
C380|Heart|967|B_Cell_Lymphomas|9679/3|Mediastinal_Large_B_cell_Lymphoma
C380|Heart|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C380|Heart|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C380|Heart|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C380|Heart|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C380|Heart|968|Diffuse_Large_B_Cell_Lymphoma|9689/3|Mucosa_associated_Lymphoma
C380|Heart|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C380|Heart|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C380|Heart|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C380|Heart|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C380|Heart|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C380|Heart|970|T_Cell_Lymphoma|9700/3|Mycosis_Fungoides
C380|Heart|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C380|Heart|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C380|Heart|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C380|Heart|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C380|Heart|970|T_Cell_Lymphoma|9709/3|Cutaneous_T_Cell_Non_Hodgkin_Lymphoma
C380|Heart|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C380|Heart|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C380|Heart|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C380|Heart|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C380|Heart|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C380|Heart|971|Adult_Non_Hodgkin_Lymphoma|9718/3|C_ALCL
C380|Heart|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C380|Heart|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C380|Heart|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C380|Heart|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C380|Heart|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C380|Heart|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C380|Heart|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C380|Heart|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C380|Heart|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C380|Heart|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C380|Heart|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C380|Heart|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C380|Heart|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C380|Heart|981|Neoplasm|9812/3|Lymphoma
C380|Heart|981|Neoplasm|9813/3|Lymphoma
C380|Heart|981|Neoplasm|9814/3|Lymphoma
C380|Heart|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C380|Heart|981|Neoplasm|9816/3|Hypodiploid_ALL
C380|Heart|981|Neoplasm|9817/3|Lymphoma
C380|Heart|981|Neoplasm|9818/3|Lymphoma
C380|Heart|981|Neoplasm|9819/3|Leukemia__B_Cell
C380|Heart|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C380|Heart|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C380|Heart|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C380|Heart|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C380|Heart|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C380|Heart|997|Neoplasm|9971/3|Polymorphic_PTLD
C380|Heart|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C381-C383, C388|Mediastinum|800|Neoplasm|8000/3|Malignant_Neoplasm
C381-C383, C388|Mediastinum|800|Neoplasm|8001/3|Malignant_Cell
C381-C383, C388|Mediastinum|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C381-C383, C388|Mediastinum|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C381-C383, C388|Mediastinum|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C381-C383, C388|Mediastinum|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C381-C383, C388|Mediastinum|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C381-C383, C388|Mediastinum|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C381-C383, C388|Mediastinum|880|Sarcoma|8800/3|Sarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C381-C383, C388|Mediastinum|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C381-C383, C388|Mediastinum|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C381-C383, C388|Mediastinum|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C381-C383, C388|Mediastinum|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C381-C383, C388|Mediastinum|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C381-C383, C388|Mediastinum|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C381-C383, C388|Mediastinum|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C381-C383, C388|Mediastinum|882|Sarcoma|8825/3|Sarcoma
C381-C383, C388|Mediastinum|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8850/3|Liposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C381-C383, C388|Mediastinum|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8855/3|Liposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C381-C383, C388|Mediastinum|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C381-C383, C388|Mediastinum|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C381-C383, C388|Mediastinum|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C381-C383, C388|Mediastinum|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C381-C383, C388|Mediastinum|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C381-C383, C388|Mediastinum|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C381-C383, C388|Mediastinum|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C381-C383, C388|Mediastinum|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C381-C383, C388|Mediastinum|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C381-C383, C388|Mediastinum|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C381-C383, C388|Mediastinum|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C381-C383, C388|Mediastinum|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C381-C383, C388|Mediastinum|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C381-C383, C388|Mediastinum|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C381-C383, C388|Mediastinum|906|Germ_Cell_Tumor|9061/3|Seminoma
C381-C383, C388|Mediastinum|906|Germ_Cell_Tumor|9062/3|Atypical_Seminoma
C381-C383, C388|Mediastinum|906|Germ_Cell_Tumor|9063/3|Testicular_Spermatocytic_Seminoma
C381-C383, C388|Mediastinum|906|Germ_Cell_Tumor|9064/3|Germinoma
C381-C383, C388|Mediastinum|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C381-C383, C388|Mediastinum|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C381-C383, C388|Mediastinum|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C381-C383, C388|Mediastinum|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C381-C383, C388|Mediastinum|908|Teratoma|9080/3|Immature_Teratoma
C381-C383, C388|Mediastinum|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C381-C383, C388|Mediastinum|908|Teratoma|9082/3|Immature_Teratoma
C381-C383, C388|Mediastinum|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C381-C383, C388|Mediastinum|908|Teratoma|9084/3|Teratoma
C381-C383, C388|Mediastinum|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C381-C383, C388|Mediastinum|910|Choriocarcinoma|9100/3|Choriocarcinoma
C381-C383, C388|Mediastinum|910|Choriocarcinoma|9101/3|Choriocarcinoma
C381-C383, C388|Mediastinum|910|Choriocarcinoma|9105/3|Epithelioid_Trophoblastic_Tumor
C381-C383, C388|Mediastinum|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9500/3|Neuroblastoma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9501/3|Medulloepithelioma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9503/3|Neuroepithelioma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C381-C383, C388|Mediastinum|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C381-C383, C388|Mediastinum|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C381-C383, C388|Mediastinum|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C381-C383, C388|Mediastinum|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C381-C383, C388|Mediastinum|957|Perineurioma|9571/3|Malignant_Perineurioma
C381-C383, C388|Mediastinum|959|Lymphoma|9590/3|Lymphoma
C381-C383, C388|Mediastinum|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C381-C383, C388|Mediastinum|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C381-C383, C388|Mediastinum|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C381-C383, C388|Mediastinum|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C381-C383, C388|Mediastinum|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C381-C383, C388|Mediastinum|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C381-C383, C388|Mediastinum|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C381-C383, C388|Mediastinum|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C381-C383, C388|Mediastinum|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C381-C383, C388|Mediastinum|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C381-C383, C388|Mediastinum|967|B_Cell_Lymphomas|9678/3|Primary_Effusion_Lymphoma
C381-C383, C388|Mediastinum|967|B_Cell_Lymphomas|9679/3|Mediastinal_Large_B_cell_Lymphoma
C381-C383, C388|Mediastinum|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C381-C383, C388|Mediastinum|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C381-C383, C388|Mediastinum|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C381-C383, C388|Mediastinum|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C381-C383, C388|Mediastinum|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C381-C383, C388|Mediastinum|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C381-C383, C388|Mediastinum|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C381-C383, C388|Mediastinum|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C381-C383, C388|Mediastinum|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C381-C383, C388|Mediastinum|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C381-C383, C388|Mediastinum|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C381-C383, C388|Mediastinum|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C381-C383, C388|Mediastinum|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C381-C383, C388|Mediastinum|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C381-C383, C388|Mediastinum|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C381-C383, C388|Mediastinum|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C381-C383, C388|Mediastinum|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C381-C383, C388|Mediastinum|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C381-C383, C388|Mediastinum|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9731/3|Plasmacytoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C381-C383, C388|Mediastinum|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C381-C383, C388|Mediastinum|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C381-C383, C388|Mediastinum|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C381-C383, C388|Mediastinum|975|Neoplasm|9750/3|Malignant_Histiocytosis
C381-C383, C388|Mediastinum|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C381-C383, C388|Mediastinum|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C381-C383, C388|Mediastinum|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C381-C383, C388|Mediastinum|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C381-C383, C388|Mediastinum|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C381-C383, C388|Mediastinum|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C381-C383, C388|Mediastinum|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C381-C383, C388|Mediastinum|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C381-C383, C388|Mediastinum|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C381-C383, C388|Mediastinum|981|Neoplasm|9812/3|Lymphoma
C381-C383, C388|Mediastinum|981|Neoplasm|9813/3|Lymphoma
C381-C383, C388|Mediastinum|981|Neoplasm|9814/3|Lymphoma
C381-C383, C388|Mediastinum|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C381-C383, C388|Mediastinum|981|Neoplasm|9816/3|Hypodiploid_ALL
C381-C383, C388|Mediastinum|981|Neoplasm|9817/3|Lymphoma
C381-C383, C388|Mediastinum|981|Neoplasm|9818/3|Lymphoma
C381-C383, C388|Mediastinum|981|Neoplasm|9819/3|Leukemia__B_Cell
C381-C383, C388|Mediastinum|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C381-C383, C388|Mediastinum|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C381-C383, C388|Mediastinum|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C381-C383, C388|Mediastinum|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C381-C383, C388|Mediastinum|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C381-C383, C388|Mediastinum|997|Neoplasm|9971/3|Polymorphic_PTLD
C381-C383, C388|Mediastinum|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C384|Pleura|800|Neoplasm|8000/3|Malignant_Neoplasm
C384|Pleura|800|Neoplasm|8001/3|Malignant_Cell
C384|Pleura|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C384|Pleura|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C384|Pleura|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C384|Pleura|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C384|Pleura|880|Sarcoma|8800/3|Sarcoma
C384|Pleura|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C384|Pleura|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C384|Pleura|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C384|Pleura|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C384|Pleura|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C384|Pleura|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C384|Pleura|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C384|Pleura|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C384|Pleura|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C384|Pleura|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C384|Pleura|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C384|Pleura|882|Sarcoma|8825/3|Sarcoma
C384|Pleura|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C384|Pleura|897|Hepatoblastoma|8973/3|Pleuropulmonary_Blastoma
C384|Pleura|905|Malignant_Mesothelioma|9050/3|Malignant_Mesothelioma
C384|Pleura|905|Malignant_Mesothelioma|9051/3|Sarcomatoid_Mesothelioma
C384|Pleura|905|Malignant_Mesothelioma|9052/3|Mesothelioma
C384|Pleura|905|Malignant_Mesothelioma|9053/3|Biphasic_Mesothelioma
C384|Pleura|959|Lymphoma|9590/3|Lymphoma
C384|Pleura|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C384|Pleura|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C384|Pleura|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C384|Pleura|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C384|Pleura|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C384|Pleura|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C384|Pleura|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C384|Pleura|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C384|Pleura|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C384|Pleura|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C384|Pleura|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C384|Pleura|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C384|Pleura|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C384|Pleura|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C384|Pleura|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C384|Pleura|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C384|Pleura|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C384|Pleura|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C384|Pleura|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C384|Pleura|967|B_Cell_Lymphomas|9678/3|Primary_Effusion_Lymphoma
C384|Pleura|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C384|Pleura|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C384|Pleura|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C384|Pleura|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C384|Pleura|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C384|Pleura|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C384|Pleura|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C384|Pleura|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C384|Pleura|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C384|Pleura|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C384|Pleura|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C384|Pleura|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C384|Pleura|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C384|Pleura|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C384|Pleura|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C384|Pleura|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C384|Pleura|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C384|Pleura|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C384|Pleura|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C384|Pleura|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C384|Pleura|973|Plasmacytoma|9731/3|Plasmacytoma
C384|Pleura|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C384|Pleura|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C384|Pleura|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C384|Pleura|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C384|Pleura|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C384|Pleura|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C384|Pleura|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C384|Pleura|975|Neoplasm|9750/3|Malignant_Histiocytosis
C384|Pleura|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C384|Pleura|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C384|Pleura|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C384|Pleura|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C384|Pleura|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C384|Pleura|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C384|Pleura|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C384|Pleura|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C384|Pleura|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C384|Pleura|981|Neoplasm|9812/3|Lymphoma
C384|Pleura|981|Neoplasm|9813/3|Lymphoma
C384|Pleura|981|Neoplasm|9814/3|Lymphoma
C384|Pleura|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C384|Pleura|981|Neoplasm|9816/3|Hypodiploid_ALL
C384|Pleura|981|Neoplasm|9817/3|Lymphoma
C384|Pleura|981|Neoplasm|9818/3|Lymphoma
C384|Pleura|981|Neoplasm|9819/3|Leukemia__B_Cell
C384|Pleura|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C384|Pleura|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C384|Pleura|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C384|Pleura|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C384|Pleura|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C384|Pleura|997|Neoplasm|9971/3|Polymorphic_PTLD
C384|Pleura|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C390,C398-C399|Respiratory_System|800|Neoplasm|8000/3|Malignant_Neoplasm
C390,C398-C399|Respiratory_System|800|Neoplasm|8001/3|Malignant_Cell
C390,C398-C399|Respiratory_System|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C390,C398-C399|Respiratory_System|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C390,C398-C399|Respiratory_System|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C390,C398-C399|Respiratory_System|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C390,C398-C399|Respiratory_System|801|Carcinoma|8010/2|In_Situ_Cancer
C390,C398-C399|Respiratory_System|801|Carcinoma|8010/3|Carcinoma
C390,C398-C399|Respiratory_System|801|Carcinoma|8011/3|Malignant_Epithelioma
C390,C398-C399|Respiratory_System|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C390,C398-C399|Respiratory_System|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C390,C398-C399|Respiratory_System|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C390,C398-C399|Respiratory_System|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C390,C398-C399|Respiratory_System|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C390,C398-C399|Respiratory_System|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C390,C398-C399|Respiratory_System|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C390,C398-C399|Respiratory_System|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C390,C398-C399|Respiratory_System|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C390,C398-C399|Respiratory_System|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C390,C398-C399|Respiratory_System|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C390,C398-C399|Respiratory_System|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C390,C398-C399|Respiratory_System|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C390,C398-C399|Respiratory_System|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C390,C398-C399|Respiratory_System|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C390,C398-C399|Respiratory_System|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C390,C398-C399|Respiratory_System|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C390,C398-C399|Respiratory_System|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C390,C398-C399|Respiratory_System|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C390,C398-C399|Respiratory_System|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C390,C398-C399|Respiratory_System|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C390,C398-C399|Respiratory_System|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C390,C398-C399|Respiratory_System|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C390,C398-C399|Respiratory_System|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C390,C398-C399|Respiratory_System|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C390,C398-C399|Respiratory_System|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C390,C398-C399|Respiratory_System|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C390,C398-C399|Respiratory_System|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C390,C398-C399|Respiratory_System|814|Adenocarcinoma|8140/3|Adenocarcinoma
C390,C398-C399|Respiratory_System|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C390,C398-C399|Respiratory_System|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C390,C398-C399|Respiratory_System|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C390,C398-C399|Respiratory_System|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C390,C398-C399|Respiratory_System|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C390,C398-C399|Respiratory_System|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C390,C398-C399|Respiratory_System|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C390,C398-C399|Respiratory_System|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C390,C398-C399|Respiratory_System|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C390,C398-C399|Respiratory_System|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C390,C398-C399|Respiratory_System|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C390,C398-C399|Respiratory_System|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C390,C398-C399|Respiratory_System|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C390,C398-C399|Respiratory_System|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C390,C398-C399|Respiratory_System|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C390,C398-C399|Respiratory_System|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C390,C398-C399|Respiratory_System|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C390,C398-C399|Respiratory_System|825|Bronchioloalveolar_Adenocarcinoma|8250/3|null
C390,C398-C399|Respiratory_System|825|Bronchioloalveolar_Adenocarcinoma|8251/3|Bronchioloalveolar_Adenocarcinoma
C390,C398-C399|Respiratory_System|825|Bronchioloalveolar_Adenocarcinoma|8252/3|Bronchioloalveolar_Adenocarcinoma
C390,C398-C399|Respiratory_System|825|Bronchioloalveolar_Adenocarcinoma|8253/3|Mucinous_Adenocarcinoma
C390,C398-C399|Respiratory_System|825|Bronchioloalveolar_Adenocarcinoma|8254/3|Adenocarcinoma
C390,C398-C399|Respiratory_System|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C390,C398-C399|Respiratory_System|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C390,C398-C399|Respiratory_System|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C390,C398-C399|Respiratory_System|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C390,C398-C399|Respiratory_System|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C390,C398-C399|Respiratory_System|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C390,C398-C399|Respiratory_System|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C390,C398-C399|Respiratory_System|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C390,C398-C399|Respiratory_System|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C390,C398-C399|Respiratory_System|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C390,C398-C399|Respiratory_System|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C390,C398-C399|Respiratory_System|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C390,C398-C399|Respiratory_System|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C390,C398-C399|Respiratory_System|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C390,C398-C399|Respiratory_System|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C390,C398-C399|Respiratory_System|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C390,C398-C399|Respiratory_System|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C390,C398-C399|Respiratory_System|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C390,C398-C399|Respiratory_System|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C390,C398-C399|Respiratory_System|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C390,C398-C399|Respiratory_System|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C390,C398-C399|Respiratory_System|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C390,C398-C399|Respiratory_System|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C390,C398-C399|Respiratory_System|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C390,C398-C399|Respiratory_System|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C390,C398-C399|Respiratory_System|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C390,C398-C399|Respiratory_System|880|Sarcoma|8800/3|Sarcoma
C390,C398-C399|Respiratory_System|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C390,C398-C399|Respiratory_System|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C390,C398-C399|Respiratory_System|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C390,C398-C399|Respiratory_System|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C390,C398-C399|Respiratory_System|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C390,C398-C399|Respiratory_System|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C390,C398-C399|Respiratory_System|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C390,C398-C399|Respiratory_System|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C390,C398-C399|Respiratory_System|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C390,C398-C399|Respiratory_System|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C390,C398-C399|Respiratory_System|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C390,C398-C399|Respiratory_System|882|Sarcoma|8825/3|Sarcoma
C390,C398-C399|Respiratory_System|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C390,C398-C399|Respiratory_System|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C390,C398-C399|Respiratory_System|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C390,C398-C399|Respiratory_System|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C390,C398-C399|Respiratory_System|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C390,C398-C399|Respiratory_System|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C390,C398-C399|Respiratory_System|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C390,C398-C399|Respiratory_System|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C390,C398-C399|Respiratory_System|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C390,C398-C399|Respiratory_System|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C390,C398-C399|Respiratory_System|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C390,C398-C399|Respiratory_System|898|Carcinosarcoma|8980/3|Carcinosarcoma
C390,C398-C399|Respiratory_System|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C390,C398-C399|Respiratory_System|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C390,C398-C399|Respiratory_System|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C390,C398-C399|Respiratory_System|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C390,C398-C399|Respiratory_System|908|Teratoma|9080/3|Immature_Teratoma
C390,C398-C399|Respiratory_System|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C390,C398-C399|Respiratory_System|908|Teratoma|9082/3|Immature_Teratoma
C390,C398-C399|Respiratory_System|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C390,C398-C399|Respiratory_System|908|Teratoma|9084/3|Teratoma
C390,C398-C399|Respiratory_System|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C390,C398-C399|Respiratory_System|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C390,C398-C399|Respiratory_System|936|Neuroepithelioma__Peripheral|9364/3|Neuroepithelioma__Peripheral
C390,C398-C399|Respiratory_System|936|Neuroepithelioma__Peripheral|9365/3|Askin_Tumor
C390,C398-C399|Respiratory_System|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|800|Neoplasm|8000/3|Malignant_Neoplasm
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|800|Neoplasm|8001/3|Malignant_Cell
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8800/3|Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|Fibromatous_Neoplasm|8812/3|Periosteal_Fibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|882|Sarcoma|8825/3|Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|884|Myxosarcoma|8840/3|Myxosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8850/3|Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8855/3|Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|904|Synovial_Sarcoma|9040/3|Synovial_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|904|Synovial_Sarcoma|9041/3|Spindle_Cell_Synovial_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|904|Synovial_Sarcoma|9042/3|Epithelial_Synovial_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|904|Synovial_Sarcoma|9043/3|Biphasic_Synovial_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9180/3|Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9181/3|Chondroblastic_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9182/3|Fibroblastic_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9183/3|Telangiectatic_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9184/3|Paget_Disease
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9185/3|Small_Cell_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9186/3|Conventional_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|918|Osteosarcoma|9187/3|Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|919|Parosteal_Osteosarcoma|9192/3|Parosteal_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|919|Parosteal_Osteosarcoma|9193/3|Periosteal_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|919|Parosteal_Osteosarcoma|9194/3|High_Grade_Surface_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|919|Parosteal_Osteosarcoma|9195/3|Conventional_Osteosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|922|Chondrosarcoma|9220/3|Chondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|922|Chondrosarcoma|9221/3|Periosteal_Chondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|923|Chondroblastoma__Malignant|9230/3|Chondroblastoma__Malignant
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|923|Chondroblastoma__Malignant|9231/3|Myxoid_Chondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|924|Neoplasm|9240/3|Mesenchymal_Chondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|924|Neoplasm|9242/3|Clear_Cell_Chondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|924|Neoplasm|9243/3|Dedifferentiated_Chondrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|925|Bone_Neoplasm|9250/3|Giant_Cell_Tumor_Of_Bone
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|925|Bone_Neoplasm|9251/3|Giant_Cell_Tumor_Of_Soft_Tissue
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|926|Ewing_Sarcoma|9260/3|Ewing_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|926|Ewing_Sarcoma|9261/3|Adamantinoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|927|Odontogenic_Neoplasm|9270/3|Malignant_Odontogenic_Tumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|929|Ameloblastic_Odontosarcoma|9290/3|Ameloblastic_Odontosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|931|Malignant_Ameloblastoma|9310/3|Malignant_Ameloblastoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|933|Ameloblastic_Fibrosarcoma|9330/3|Ameloblastic_Fibrosarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|934|Malignant_Odontogenic_Tumor|9342/3|Malignant_Odontogenic_Tumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|936|Neuroepithelioma__Peripheral|9364/3|Neuroepithelioma__Peripheral
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|936|Neuroepithelioma__Peripheral|9365/3|Askin_Tumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|937|Chordoma|9370/3|Chordoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|937|Chordoma|9371/3|Chondroid_Chordoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|959|Lymphoma|9590/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9731/3|Plasmacytoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9732/3|Plasma_Cell_Myeloma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|Neoplasm|9750/3|Malignant_Histiocytosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9812/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9813/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9814/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9816/3|Hypodiploid_ALL
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9817/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9818/3|Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|981|Neoplasm|9819/3|Leukemia__B_Cell
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|997|Neoplasm|9971/3|Polymorphic_PTLD
C400-C403,C408-C409,C412-C414,C418-C419|Mandible|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C410|Skull|800|Neoplasm|8000/3|Malignant_Neoplasm
C410|Skull|800|Neoplasm|8001/3|Malignant_Cell
C410|Skull|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C410|Skull|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C410|Skull|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C410|Skull|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C410|Skull|880|Sarcoma|8800/3|Sarcoma
C410|Skull|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C410|Skull|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C410|Skull|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C410|Skull|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C410|Skull|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C410|Skull|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C410|Skull|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C410|Skull|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C410|Skull|881|Fibromatous_Neoplasm|8812/3|Periosteal_Fibrosarcoma
C410|Skull|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C410|Skull|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C410|Skull|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C410|Skull|882|Sarcoma|8825/3|Sarcoma
C410|Skull|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C410|Skull|884|Myxosarcoma|8840/3|Myxosarcoma
C410|Skull|885|Liposarcoma|8850/3|Liposarcoma
C410|Skull|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C410|Skull|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C410|Skull|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C410|Skull|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C410|Skull|885|Liposarcoma|8855/3|Liposarcoma
C410|Skull|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C410|Skull|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C410|Skull|904|Synovial_Sarcoma|9040/3|Synovial_Sarcoma
C410|Skull|904|Synovial_Sarcoma|9041/3|Spindle_Cell_Synovial_Sarcoma
C410|Skull|904|Synovial_Sarcoma|9042/3|Epithelial_Synovial_Sarcoma
C410|Skull|904|Synovial_Sarcoma|9043/3|Biphasic_Synovial_Sarcoma
C410|Skull|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C410|Skull|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C410|Skull|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C410|Skull|918|Osteosarcoma|9180/3|Osteosarcoma
C410|Skull|918|Osteosarcoma|9181/3|Chondroblastic_Osteosarcoma
C410|Skull|918|Osteosarcoma|9182/3|Fibroblastic_Osteosarcoma
C410|Skull|918|Osteosarcoma|9183/3|Telangiectatic_Osteosarcoma
C410|Skull|918|Osteosarcoma|9184/3|Paget_Disease
C410|Skull|918|Osteosarcoma|9185/3|Small_Cell_Osteosarcoma
C410|Skull|918|Osteosarcoma|9186/3|Conventional_Osteosarcoma
C410|Skull|918|Osteosarcoma|9187/3|Osteosarcoma
C410|Skull|919|Parosteal_Osteosarcoma|9192/3|Parosteal_Osteosarcoma
C410|Skull|919|Parosteal_Osteosarcoma|9193/3|Periosteal_Osteosarcoma
C410|Skull|919|Parosteal_Osteosarcoma|9194/3|High_Grade_Surface_Osteosarcoma
C410|Skull|919|Parosteal_Osteosarcoma|9195/3|Conventional_Osteosarcoma
C410|Skull|922|Chondrosarcoma|9220/3|Chondrosarcoma
C410|Skull|922|Chondrosarcoma|9221/3|Periosteal_Chondrosarcoma
C410|Skull|923|Chondroblastoma__Malignant|9230/3|Chondroblastoma__Malignant
C410|Skull|923|Chondroblastoma__Malignant|9231/3|Myxoid_Chondrosarcoma
C410|Skull|924|Neoplasm|9240/3|Mesenchymal_Chondrosarcoma
C410|Skull|924|Neoplasm|9242/3|Clear_Cell_Chondrosarcoma
C410|Skull|924|Neoplasm|9243/3|Dedifferentiated_Chondrosarcoma
C410|Skull|925|Bone_Neoplasm|9250/3|Giant_Cell_Tumor_Of_Bone
C410|Skull|925|Bone_Neoplasm|9251/3|Giant_Cell_Tumor_Of_Soft_Tissue
C410|Skull|926|Ewing_Sarcoma|9260/3|Ewing_Sarcoma
C410|Skull|926|Ewing_Sarcoma|9261/3|Adamantinoma
C410|Skull|927|Odontogenic_Neoplasm|9270/3|Malignant_Odontogenic_Tumor
C410|Skull|929|Ameloblastic_Odontosarcoma|9290/3|Ameloblastic_Odontosarcoma
C410|Skull|930|Odontogenic_Neoplasm|9302/3|Ghost_Cell_Odontogenic_Carcinoma
C410|Skull|931|Malignant_Ameloblastoma|9310/3|Malignant_Ameloblastoma
C410|Skull|933|Ameloblastic_Fibrosarcoma|9330/3|Ameloblastic_Fibrosarcoma
C410|Skull|934|Malignant_Odontogenic_Tumor|9341/3|Clear_Cell_Odontogenic_Carcinoma
C410|Skull|934|Malignant_Odontogenic_Tumor|9342/3|Malignant_Odontogenic_Tumor
C410|Skull|936|Neuroepithelioma__Peripheral|9364/3|Neuroepithelioma__Peripheral
C410|Skull|936|Neuroepithelioma__Peripheral|9365/3|Askin_Tumor
C410|Skull|937|Chordoma|9370/3|Chordoma
C410|Skull|937|Chordoma|9371/3|Chondroid_Chordoma
C410|Skull|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C410|Skull|959|Lymphoma|9590/3|Lymphoma
C410|Skull|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C410|Skull|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C410|Skull|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C410|Skull|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C410|Skull|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C410|Skull|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C410|Skull|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C410|Skull|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C410|Skull|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C410|Skull|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C410|Skull|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C410|Skull|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C410|Skull|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C410|Skull|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C410|Skull|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C410|Skull|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C410|Skull|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C410|Skull|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C410|Skull|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C410|Skull|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C410|Skull|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C410|Skull|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C410|Skull|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C410|Skull|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C410|Skull|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C410|Skull|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C410|Skull|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C410|Skull|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C410|Skull|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C410|Skull|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C410|Skull|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C410|Skull|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C410|Skull|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C410|Skull|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C410|Skull|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C410|Skull|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C410|Skull|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C410|Skull|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C410|Skull|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C410|Skull|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C410|Skull|973|Plasmacytoma|9731/3|Plasmacytoma
C410|Skull|973|Plasmacytoma|9732/3|Plasma_Cell_Myeloma
C410|Skull|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C410|Skull|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C410|Skull|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C410|Skull|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C410|Skull|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C410|Skull|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C410|Skull|975|Neoplasm|9750/3|Malignant_Histiocytosis
C410|Skull|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C410|Skull|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C410|Skull|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C410|Skull|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C410|Skull|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C410|Skull|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C410|Skull|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C410|Skull|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C410|Skull|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C410|Skull|981|Neoplasm|9812/3|Lymphoma
C410|Skull|981|Neoplasm|9813/3|Lymphoma
C410|Skull|981|Neoplasm|9814/3|Lymphoma
C410|Skull|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C410|Skull|981|Neoplasm|9816/3|Hypodiploid_ALL
C410|Skull|981|Neoplasm|9817/3|Lymphoma
C410|Skull|981|Neoplasm|9818/3|Lymphoma
C410|Skull|981|Neoplasm|9819/3|Leukemia__B_Cell
C410|Skull|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C410|Skull|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C410|Skull|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C410|Skull|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C410|Skull|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C410|Skull|997|Neoplasm|9971/3|Polymorphic_PTLD
C410|Skull|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C411|Mandible|800|Neoplasm|8000/3|Malignant_Neoplasm
C411|Mandible|800|Neoplasm|8001/3|Malignant_Cell
C411|Mandible|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C411|Mandible|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C411|Mandible|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C411|Mandible|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C411|Mandible|880|Sarcoma|8800/3|Sarcoma
C411|Mandible|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C411|Mandible|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C411|Mandible|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C411|Mandible|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C411|Mandible|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C411|Mandible|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C411|Mandible|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C411|Mandible|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C411|Mandible|881|Fibromatous_Neoplasm|8812/3|Periosteal_Fibrosarcoma
C411|Mandible|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C411|Mandible|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C411|Mandible|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C411|Mandible|882|Sarcoma|8825/3|Sarcoma
C411|Mandible|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C411|Mandible|884|Myxosarcoma|8840/3|Myxosarcoma
C411|Mandible|885|Liposarcoma|8850/3|Liposarcoma
C411|Mandible|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C411|Mandible|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C411|Mandible|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C411|Mandible|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C411|Mandible|885|Liposarcoma|8855/3|Liposarcoma
C411|Mandible|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C411|Mandible|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C411|Mandible|904|Synovial_Sarcoma|9040/3|Synovial_Sarcoma
C411|Mandible|904|Synovial_Sarcoma|9041/3|Spindle_Cell_Synovial_Sarcoma
C411|Mandible|904|Synovial_Sarcoma|9042/3|Epithelial_Synovial_Sarcoma
C411|Mandible|904|Synovial_Sarcoma|9043/3|Biphasic_Synovial_Sarcoma
C411|Mandible|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C411|Mandible|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C411|Mandible|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C411|Mandible|918|Osteosarcoma|9180/3|Osteosarcoma
C411|Mandible|918|Osteosarcoma|9181/3|Chondroblastic_Osteosarcoma
C411|Mandible|918|Osteosarcoma|9182/3|Fibroblastic_Osteosarcoma
C411|Mandible|918|Osteosarcoma|9183/3|Telangiectatic_Osteosarcoma
C411|Mandible|918|Osteosarcoma|9184/3|Paget_Disease
C411|Mandible|918|Osteosarcoma|9185/3|Small_Cell_Osteosarcoma
C411|Mandible|918|Osteosarcoma|9186/3|Conventional_Osteosarcoma
C411|Mandible|918|Osteosarcoma|9187/3|Osteosarcoma
C411|Mandible|919|Parosteal_Osteosarcoma|9192/3|Parosteal_Osteosarcoma
C411|Mandible|919|Parosteal_Osteosarcoma|9193/3|Periosteal_Osteosarcoma
C411|Mandible|919|Parosteal_Osteosarcoma|9194/3|High_Grade_Surface_Osteosarcoma
C411|Mandible|919|Parosteal_Osteosarcoma|9195/3|Conventional_Osteosarcoma
C411|Mandible|922|Chondrosarcoma|9220/3|Chondrosarcoma
C411|Mandible|922|Chondrosarcoma|9221/3|Periosteal_Chondrosarcoma
C411|Mandible|923|Chondroblastoma__Malignant|9230/3|Chondroblastoma__Malignant
C411|Mandible|923|Chondroblastoma__Malignant|9231/3|Myxoid_Chondrosarcoma
C411|Mandible|924|Neoplasm|9240/3|Mesenchymal_Chondrosarcoma
C411|Mandible|924|Neoplasm|9242/3|Clear_Cell_Chondrosarcoma
C411|Mandible|924|Neoplasm|9243/3|Dedifferentiated_Chondrosarcoma
C411|Mandible|925|Bone_Neoplasm|9250/3|Giant_Cell_Tumor_Of_Bone
C411|Mandible|925|Bone_Neoplasm|9251/3|Giant_Cell_Tumor_Of_Soft_Tissue
C411|Mandible|926|Ewing_Sarcoma|9260/3|Ewing_Sarcoma
C411|Mandible|926|Ewing_Sarcoma|9261/3|Adamantinoma
C411|Mandible|927|Odontogenic_Neoplasm|9270/3|Malignant_Odontogenic_Tumor
C411|Mandible|929|Ameloblastic_Odontosarcoma|9290/3|Ameloblastic_Odontosarcoma
C411|Mandible|930|Odontogenic_Neoplasm|9302/3|Ghost_Cell_Odontogenic_Carcinoma
C411|Mandible|931|Malignant_Ameloblastoma|9310/3|Malignant_Ameloblastoma
C411|Mandible|933|Ameloblastic_Fibrosarcoma|9330/3|Ameloblastic_Fibrosarcoma
C411|Mandible|934|Malignant_Odontogenic_Tumor|9341/3|Clear_Cell_Odontogenic_Carcinoma
C411|Mandible|934|Malignant_Odontogenic_Tumor|9342/3|Malignant_Odontogenic_Tumor
C411|Mandible|936|Neuroepithelioma__Peripheral|9364/3|Neuroepithelioma__Peripheral
C411|Mandible|936|Neuroepithelioma__Peripheral|9365/3|Askin_Tumor
C411|Mandible|937|Chordoma|9370/3|Chordoma
C411|Mandible|937|Chordoma|9371/3|Chondroid_Chordoma
C411|Mandible|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C411|Mandible|959|Lymphoma|9590/3|Lymphoma
C411|Mandible|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C411|Mandible|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C411|Mandible|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C411|Mandible|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C411|Mandible|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C411|Mandible|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C411|Mandible|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C411|Mandible|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C411|Mandible|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C411|Mandible|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C411|Mandible|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C411|Mandible|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C411|Mandible|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C411|Mandible|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C411|Mandible|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C411|Mandible|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C411|Mandible|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C411|Mandible|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C411|Mandible|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C411|Mandible|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C411|Mandible|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C411|Mandible|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C411|Mandible|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C411|Mandible|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C411|Mandible|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C411|Mandible|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C411|Mandible|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C411|Mandible|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C411|Mandible|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C411|Mandible|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C411|Mandible|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C411|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C411|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C411|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C411|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C411|Mandible|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C411|Mandible|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C411|Mandible|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C411|Mandible|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C411|Mandible|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C411|Mandible|973|Plasmacytoma|9731/3|Plasmacytoma
C411|Mandible|973|Plasmacytoma|9732/3|Plasma_Cell_Myeloma
C411|Mandible|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C411|Mandible|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C411|Mandible|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C411|Mandible|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C411|Mandible|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C411|Mandible|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C411|Mandible|975|Neoplasm|9750/3|Malignant_Histiocytosis
C411|Mandible|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C411|Mandible|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C411|Mandible|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C411|Mandible|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C411|Mandible|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C411|Mandible|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C411|Mandible|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C411|Mandible|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C411|Mandible|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C411|Mandible|981|Neoplasm|9812/3|Lymphoma
C411|Mandible|981|Neoplasm|9813/3|Lymphoma
C411|Mandible|981|Neoplasm|9814/3|Lymphoma
C411|Mandible|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C411|Mandible|981|Neoplasm|9816/3|Hypodiploid_ALL
C411|Mandible|981|Neoplasm|9817/3|Lymphoma
C411|Mandible|981|Neoplasm|9818/3|Lymphoma
C411|Mandible|981|Neoplasm|9819/3|Leukemia__B_Cell
C411|Mandible|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C411|Mandible|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C411|Mandible|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C411|Mandible|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C411|Mandible|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C411|Mandible|997|Neoplasm|9971/3|Polymorphic_PTLD
C411|Mandible|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C420, C421, C424|Bone_Marrow|959|Lymphoma|9590/3|Lymphoma
C420, C421, C424|Bone_Marrow|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C420, C421, C424|Bone_Marrow|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C420, C421, C424|Bone_Marrow|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C420, C421, C424|Bone_Marrow|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C420, C421, C424|Bone_Marrow|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C420, C421, C424|Bone_Marrow|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C420, C421, C424|Bone_Marrow|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C420, C421, C424|Bone_Marrow|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C420, C421, C424|Bone_Marrow|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C420, C421, C424|Bone_Marrow|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C420, C421, C424|Bone_Marrow|967|B_Cell_Lymphomas|9678/3|Primary_Effusion_Lymphoma
C420, C421, C424|Bone_Marrow|967|B_Cell_Lymphomas|9679/3|Mediastinal_Large_B_cell_Lymphoma
C420, C421, C424|Bone_Marrow|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C420, C421, C424|Bone_Marrow|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C420, C421, C424|Bone_Marrow|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C420, C421, C424|Bone_Marrow|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|968|Diffuse_Large_B_Cell_Lymphoma|9689/3|Mucosa_associated_Lymphoma
C420, C421, C424|Bone_Marrow|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C420, C421, C424|Bone_Marrow|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C420, C421, C424|Bone_Marrow|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C420, C421, C424|Bone_Marrow|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C420, C421, C424|Bone_Marrow|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C420, C421, C424|Bone_Marrow|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C420, C421, C424|Bone_Marrow|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C420, C421, C424|Bone_Marrow|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C420, C421, C424|Bone_Marrow|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C420, C421, C424|Bone_Marrow|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C420, C421, C424|Bone_Marrow|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C420, C421, C424|Bone_Marrow|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C420, C421, C424|Bone_Marrow|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C420, C421, C424|Bone_Marrow|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C420, C421, C424|Bone_Marrow|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C420, C421, C424|Bone_Marrow|973|Plasmacytoma|9731/3|Plasmacytoma
C420, C421, C424|Bone_Marrow|973|Plasmacytoma|9732/3|Plasma_Cell_Myeloma
C420, C421, C424|Bone_Marrow|973|Plasmacytoma|9733/3|Plasma_Cell_Leukemia
C420, C421, C424|Bone_Marrow|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C420, C421, C424|Bone_Marrow|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C420, C421, C424|Bone_Marrow|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C420, C421, C424|Bone_Marrow|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C420, C421, C424|Bone_Marrow|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C420, C421, C424|Bone_Marrow|974|Mast_Cell_Neoplasm|9742/3|Mast_Cell_Leukemia
C420, C421, C424|Bone_Marrow|975|Neoplasm|9750/3|Malignant_Histiocytosis
C420, C421, C424|Bone_Marrow|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C420, C421, C424|Bone_Marrow|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C420, C421, C424|Bone_Marrow|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C420, C421, C424|Bone_Marrow|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C420, C421, C424|Bone_Marrow|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C420, C421, C424|Bone_Marrow|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C420, C421, C424|Bone_Marrow|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C420, C421, C424|Bone_Marrow|976|Immunoproliferative_Disorder|9760/3|Immunoproliferative_Disorder
C420, C421, C424|Bone_Marrow|976|Immunoproliferative_Disorder|9761/3|Waldenstrom_Macroglobulinemia
C420, C421, C424|Bone_Marrow|976|Immunoproliferative_Disorder|9762/3|Heavy_Chain_Disease
C420, C421, C424|Bone_Marrow|980|Leukemia|9800/3|Leukemia
C420, C421, C424|Bone_Marrow|980|Leukemia|9801/3|Acute_Leukemia
C420, C421, C424|Bone_Marrow|980|Leukemia|9805/3|Acute_Biphenotypic_Leukemia
C420, C421, C424|Bone_Marrow|980|Leukemia|9806/3|Mixed_Phenotype_Acute_Leukemia
C420, C421, C424|Bone_Marrow|980|Leukemia|9807/3|Mixed_Phenotype_Acute_Leukemia
C420, C421, C424|Bone_Marrow|980|Leukemia|9808/3|Mixed_Phenotype_Acute_Leukemia
C420, C421, C424|Bone_Marrow|980|Leukemia|9809/3|Mixed_Phenotype_Acute_Leukemia
C420, C421, C424|Bone_Marrow|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C420, C421, C424|Bone_Marrow|981|Neoplasm|9812/3|Lymphoma
C420, C421, C424|Bone_Marrow|981|Neoplasm|9813/3|Lymphoma
C420, C421, C424|Bone_Marrow|981|Neoplasm|9814/3|Lymphoma
C420, C421, C424|Bone_Marrow|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C420, C421, C424|Bone_Marrow|981|Neoplasm|9816/3|Hypodiploid_ALL
C420, C421, C424|Bone_Marrow|981|Neoplasm|9817/3|Lymphoma
C420, C421, C424|Bone_Marrow|981|Neoplasm|9818/3|Lymphoma
C420, C421, C424|Bone_Marrow|981|Neoplasm|9819/3|Leukemia__B_Cell
C420, C421, C424|Bone_Marrow|982|Lymphoid_Leukemia|9820/3|Lymphoid_Leukemia
C420, C421, C424|Bone_Marrow|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C420, C421, C424|Bone_Marrow|982|Lymphoid_Leukemia|9826/3|Burkitt_Leukemia
C420, C421, C424|Bone_Marrow|982|Lymphoid_Leukemia|9827/3|Adult_T_cell_Leukemia
C420, C421, C424|Bone_Marrow|982|Lymphoid_Leukemia|9828/3|L2_Acute_Lymphoblastic_Leukemia
C420, C421, C424|Bone_Marrow|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C420, C421, C424|Bone_Marrow|983|Leukemia|9832/3|Prolymphocytic_Leukemia
C420, C421, C424|Bone_Marrow|983|Leukemia|9833/3|B_Cell_Prolymphocytic_Leukemia
C420, C421, C424|Bone_Marrow|983|Leukemia|9834/3|T_Cell_Prolymphocytic_Leukemia
C420, C421, C424|Bone_Marrow|983|Leukemia|9835/3|Acute_Lymphoblastic_Leukemia
C420, C421, C424|Bone_Marrow|983|Leukemia|9836/3|B_Acute_Lymphoblastic_Leukemia
C420, C421, C424|Bone_Marrow|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C420, C421, C424|Bone_Marrow|984|Leukemia|9840/3|Acute_Erythroid_Leukemia
C420, C421, C424|Bone_Marrow|986|Myeloid_Leukemia|9860/3|Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|986|Myeloid_Leukemia|9861/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|986|Myeloid_Leukemia|9863/3|Myeloid_Leukemia__Chronic
C420, C421, C424|Bone_Marrow|986|Myeloid_Leukemia|9865/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|986|Myeloid_Leukemia|9866/3|Acute_Promyelocytic_Leukemia
C420, C421, C424|Bone_Marrow|986|Myeloid_Leukemia|9867/3|Acute_Myelomonocytic_Leukemia
C420, C421, C424|Bone_Marrow|986|Myeloid_Leukemia|9869/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9870/3|Acute_Basophilic_Leukemia
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9871/3|CMML_With_Eosinophilia
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9872/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9873/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9874/3|Acute_Myeloid_Leukemia_With_Maturation
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9875/3|Myeloid_Leukemia__Chronic
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9876/3|Subacute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9877/3|Acute_Myeloid_Leukemia_With_Mutated_NPM1
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9878/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|987|Myeloid_Leukemia|9879/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|989|Leukemia|9891/3|Acute_Monocytic_Leukemia
C420, C421, C424|Bone_Marrow|989|Leukemia|9895/3|AML_With_Multilineage_Dysplasia
C420, C421, C424|Bone_Marrow|989|Leukemia|9896/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|989|Leukemia|9897/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|989|Leukemia|9898/3|Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|991|Acute_Megakaryocytic_Leukemias|9910/3|Acute_Megakaryocytic_Leukemias
C420, C421, C424|Bone_Marrow|991|Acute_Megakaryocytic_Leukemias|9911/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|991|Acute_Megakaryocytic_Leukemias|9912/3|Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|992|Therapy_Related_Leukemia|9920/3|Therapy_Related_Acute_Myeloid_Leukemia
C420, C421, C424|Bone_Marrow|993|Myeloid_Sarcoma|9930/3|Myeloid_Sarcoma
C420, C421, C424|Bone_Marrow|993|Myeloid_Sarcoma|9931/3|Acute_Panmyelosis_With_Myelofibrosis
C420, C421, C424|Bone_Marrow|994|Leukemia|9940/3|Hairy_Cell_Leukemia
C420, C421, C424|Bone_Marrow|994|Leukemia|9945/3|Chronic_Myelomonocytic_Leukemia
C420, C421, C424|Bone_Marrow|994|Leukemia|9946/3|Juvenile_Myelomonocytic_Leukemia
C420, C421, C424|Bone_Marrow|994|Leukemia|9948/3|Aggressive_NK_Cell_Leukemia
C420, C421, C424|Bone_Marrow|995|Polycythemia_Vera|9950/3|Polycythemia_Vera
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9960/3|Myeloproliferative_Neoplasm
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9961/3|Primary_Myelofibrosis
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9962/3|Essential_Thrombocythemia
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9963/3|Chronic_Neutrophilic_Leukemia
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9964/3|Hypereosinophilic_Syndrome
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9966/3|Neoplasm
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C420, C421, C424|Bone_Marrow|996|Myeloproliferative_Neoplasm|9968/3|Lymphocytic_Neoplasm
C420, C421, C424|Bone_Marrow|997|Neoplasm|9971/3|Polymorphic_PTLD
C420, C421, C424|Bone_Marrow|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C420, C421, C424|Bone_Marrow|998|Refractory_Anemia|9980/3|Refractory_Anemia
C420, C421, C424|Bone_Marrow|998|Refractory_Anemia|9982/3|Refractory_Anemia_With_Sideroblasts
C420, C421, C424|Bone_Marrow|998|Refractory_Anemia|9983/3|Refractory_Anemia_With_Excess_Blasts
C420, C421, C424|Bone_Marrow|998|Refractory_Anemia|9984/3|Refractory_Anemia_With_Excess_Blasts
C420, C421, C424|Bone_Marrow|998|Refractory_Anemia|9985/3|Refractory_Cytopenia_Of_Childhood
C420, C421, C424|Bone_Marrow|998|Refractory_Anemia|9986/3|_5q_syndrome
C420, C421, C424|Bone_Marrow|998|Refractory_Anemia|9987/3|Myelodysplastic_Syndrome
C420, C421, C424|Bone_Marrow|998|Refractory_Anemia|9989/3|Myelodysplastic_Syndrome
C420, C421, C424|Bone_Marrow|999|Myelodysplastic_Syndrome|9991/3|Refractory_Neutropenia
C420, C421, C424|Bone_Marrow|999|Myelodysplastic_Syndrome|9992/3|Refractory_Thrombocytopenia
C420, C421, C424|Bone_Marrow|999|Myelodysplastic_Syndrome|9993/3|Myelodysplastic_Syndrome
C422|Spleen|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C422|Spleen|959|Lymphoma|9590/3|Lymphoma
C422|Spleen|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C422|Spleen|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C422|Spleen|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C422|Spleen|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C422|Spleen|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C422|Spleen|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C422|Spleen|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C422|Spleen|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C422|Spleen|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C422|Spleen|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C422|Spleen|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C422|Spleen|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C422|Spleen|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C422|Spleen|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C422|Spleen|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C422|Spleen|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C422|Spleen|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C422|Spleen|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C422|Spleen|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C422|Spleen|967|B_Cell_Lymphomas|9678/3|Primary_Effusion_Lymphoma
C422|Spleen|967|B_Cell_Lymphomas|9679/3|Mediastinal_Large_B_cell_Lymphoma
C422|Spleen|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C422|Spleen|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C422|Spleen|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C422|Spleen|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C422|Spleen|968|Diffuse_Large_B_Cell_Lymphoma|9689/3|Mucosa_associated_Lymphoma
C422|Spleen|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C422|Spleen|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C422|Spleen|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C422|Spleen|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C422|Spleen|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C422|Spleen|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C422|Spleen|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C422|Spleen|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C422|Spleen|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C422|Spleen|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C422|Spleen|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C422|Spleen|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C422|Spleen|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C422|Spleen|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C422|Spleen|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C422|Spleen|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C422|Spleen|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C422|Spleen|973|Plasmacytoma|9731/3|Plasmacytoma
C422|Spleen|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C422|Spleen|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C422|Spleen|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C422|Spleen|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C422|Spleen|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C422|Spleen|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C422|Spleen|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C422|Spleen|975|Neoplasm|9750/3|Malignant_Histiocytosis
C422|Spleen|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C422|Spleen|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C422|Spleen|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C422|Spleen|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C422|Spleen|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C422|Spleen|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C422|Spleen|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C422|Spleen|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C422|Spleen|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C422|Spleen|981|Neoplasm|9812/3|Lymphoma
C422|Spleen|981|Neoplasm|9813/3|Lymphoma
C422|Spleen|981|Neoplasm|9814/3|Lymphoma
C422|Spleen|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C422|Spleen|981|Neoplasm|9816/3|Hypodiploid_ALL
C422|Spleen|981|Neoplasm|9817/3|Lymphoma
C422|Spleen|981|Neoplasm|9818/3|Lymphoma
C422|Spleen|981|Neoplasm|9819/3|Leukemia__B_Cell
C422|Spleen|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C422|Spleen|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C422|Spleen|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C422|Spleen|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C422|Spleen|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C422|Spleen|997|Neoplasm|9971/3|Polymorphic_PTLD
C422|Spleen|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C423|Reticuloendothelial_System|959|Lymphoma|9590/3|Lymphoma
C423|Reticuloendothelial_System|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C423|Reticuloendothelial_System|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C423|Reticuloendothelial_System|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C423|Reticuloendothelial_System|975|Neoplasm|9750/3|Malignant_Histiocytosis
C423|Reticuloendothelial_System|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C423|Reticuloendothelial_System|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C423|Reticuloendothelial_System|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C423|Reticuloendothelial_System|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C423|Reticuloendothelial_System|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C423|Reticuloendothelial_System|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C440-C449|Skin|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C440-C449|Skin|811|Pilomatrical_Carcinoma|8110/3|Pilomatrical_Carcinoma
C440-C449|Skin|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C440-C449|Skin|814|Adenocarcinoma|8140/3|Adenocarcinoma
C440-C449|Skin|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C440-C449|Skin|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C440-C449|Skin|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C440-C449|Skin|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C440-C449|Skin|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C440-C449|Skin|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C440-C449|Skin|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C440-C449|Skin|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C440-C449|Skin|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C440-C449|Skin|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C440-C449|Skin|824|Atypical_Carcinoid_Tumor|8247/3|Merkel_Cell_Carcinoma
C440-C449|Skin|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C440-C449|Skin|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C440-C449|Skin|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C440-C449|Skin|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C440-C449|Skin|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C440-C449|Skin|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C440-C449|Skin|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C440-C449|Skin|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C440-C449|Skin|839|Adnexal_Carcinoma|8390/3|Adnexal_Carcinoma
C440-C449|Skin|840|Sweat_Gland_Adenocarcinoma|8400/3|Sweat_Gland_Adenocarcinoma
C440-C449|Skin|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C440-C449|Skin|840|Sweat_Gland_Adenocarcinoma|8402/3|Sweat_Gland_Adenocarcinoma
C440-C449|Skin|840|Sweat_Gland_Adenocarcinoma|8403/3|Spiradenocarcinoma
C440-C449|Skin|840|Sweat_Gland_Adenocarcinoma|8407/3|Microcystic_Adnexal_Carcinoma
C440-C449|Skin|840|Sweat_Gland_Adenocarcinoma|8408/3|Digital_Papillary_Eccrine_Carcinoma
C440-C449|Skin|840|Sweat_Gland_Adenocarcinoma|8409/3|Eccrine_Porocarcinoma
C440-C449|Skin|841|Eccrine_Adenocarcinoma|8410/3|Sebaceous_Adenocarcinoma
C440-C449|Skin|841|Eccrine_Adenocarcinoma|8413/3|Eccrine_Adenocarcinoma
C440-C449|Skin|842|Ceruminous_Adenocarcinoma|8420/3|Ceruminous_Adenocarcinoma
C440-C449|Skin|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C440-C449|Skin|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C440-C449|Skin|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C440-C449|Skin|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C440-C449|Skin|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C440-C449|Skin|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C440-C449|Skin|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C440-C449|Skin|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C440-C449|Skin|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C440-C449|Skin|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C440-C449|Skin|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C440-C449|Skin|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C440-C449|Skin|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C440-C449|Skin|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C440-C449|Skin|872|Melanoma|8720/3|Melanoma
C440-C449|Skin|872|Melanoma|8721/3|Nodular_Melanoma
C440-C449|Skin|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C440-C449|Skin|872|Melanoma|8723/3|Regressing_Melanoma
C440-C449|Skin|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C440-C449|Skin|874|Nevus|8740/3|Melanoma_In_Junctional_Nevus
C440-C449|Skin|874|Nevus|8741/2|Precancerous_Melanosis
C440-C449|Skin|874|Nevus|8741/3|Melanoma
C440-C449|Skin|874|Nevus|8742/2|Lentigo_Maligna
C440-C449|Skin|874|Nevus|8742/3|Lentigo_Maligna_Melanoma
C440-C449|Skin|874|Nevus|8743/2|Superficial_Spreading_Melanoma
C440-C449|Skin|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C440-C449|Skin|874|Nevus|8744/3|Acral_Lentiginous_Melanoma
C440-C449|Skin|874|Nevus|8745/3|Desmoplastic_Melanoma
C440-C449|Skin|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C440-C449|Skin|876|Nevus|8761/3|Giant_Congenital_Nevus
C440-C449|Skin|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C440-C449|Skin|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C440-C449|Skin|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C440-C449|Skin|878|Melanoma_Arising_From_Blue_Nevus|8780/3|Melanoma_Arising_From_Blue_Nevus
C440-C449|Skin|880|Sarcoma|8800/3|Sarcoma
C440-C449|Skin|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C440-C449|Skin|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C440-C449|Skin|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C440-C449|Skin|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C440-C449|Skin|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C440-C449|Skin|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C440-C449|Skin|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C440-C449|Skin|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C440-C449|Skin|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C440-C449|Skin|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C440-C449|Skin|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C440-C449|Skin|882|Sarcoma|8825/3|Sarcoma
C440-C449|Skin|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C440-C449|Skin|883|Benign_Fibrous_Histiocytoma|8832/3|Dermatofibrosarcoma_Protuberans
C440-C449|Skin|883|Benign_Fibrous_Histiocytoma|8833/3|Dermatofibrosarcoma_Protuberans
C440-C449|Skin|885|Liposarcoma|8850/3|Liposarcoma
C440-C449|Skin|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C440-C449|Skin|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C440-C449|Skin|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C440-C449|Skin|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C440-C449|Skin|885|Liposarcoma|8855/3|Liposarcoma
C440-C449|Skin|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C440-C449|Skin|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C440-C449|Skin|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C440-C449|Skin|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C440-C449|Skin|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C440-C449|Skin|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C440-C449|Skin|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C440-C449|Skin|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C440-C449|Skin|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C440-C449|Skin|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C440-C449|Skin|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C440-C449|Skin|898|Carcinosarcoma|8980/3|Carcinosarcoma
C440-C449|Skin|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C440-C449|Skin|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C440-C449|Skin|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C440-C449|Skin|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C440-C449|Skin|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C440-C449|Skin|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C440-C449|Skin|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C440-C449|Skin|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C440-C449|Skin|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C440-C449|Skin|959|Lymphoma|9590/3|Lymphoma
C440-C449|Skin|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C440-C449|Skin|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C440-C449|Skin|959|Lymphoma|9597/3|Crosti_s_Disease
C440-C449|Skin|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C440-C449|Skin|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C440-C449|Skin|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C440-C449|Skin|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C440-C449|Skin|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C440-C449|Skin|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C440-C449|Skin|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C440-C449|Skin|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C440-C449|Skin|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C440-C449|Skin|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C440-C449|Skin|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C440-C449|Skin|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C440-C449|Skin|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C440-C449|Skin|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C440-C449|Skin|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C440-C449|Skin|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C440-C449|Skin|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C440-C449|Skin|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C440-C449|Skin|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C440-C449|Skin|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C440-C449|Skin|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C440-C449|Skin|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C440-C449|Skin|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C440-C449|Skin|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C440-C449|Skin|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C440-C449|Skin|970|T_Cell_Lymphoma|9700/3|Mycosis_Fungoides
C440-C449|Skin|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C440-C449|Skin|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C440-C449|Skin|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C440-C449|Skin|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C440-C449|Skin|970|T_Cell_Lymphoma|9709/3|Cutaneous_T_Cell_Non_Hodgkin_Lymphoma
C440-C449|Skin|971|Adult_Non_Hodgkin_Lymphoma|9718/3|C_ALCL
C440-C449|Skin|972|Lymphoblastic_Lymphoma|9725/3|Hydroa_Vacciniforme_Like_Lymphoma
C440-C449|Skin|972|Lymphoblastic_Lymphoma|9726/3|T_Cell_Lymphoma
C440-C449|Skin|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C440-C449|Skin|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C440-C449|Skin|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C440-C449|Skin|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C440-C449|Skin|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C440-C449|Skin|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|800|Neoplasm|8000/3|Malignant_Neoplasm
C470-C476,C478-C479|Peripheral_Nerve|800|Neoplasm|8001/3|Malignant_Cell
C470-C476,C478-C479|Peripheral_Nerve|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C470-C476,C478-C479|Peripheral_Nerve|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C470-C476,C478-C479|Peripheral_Nerve|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C470-C476,C478-C479|Peripheral_Nerve|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C470-C476,C478-C479|Peripheral_Nerve|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C470-C476,C478-C479|Peripheral_Nerve|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C470-C476,C478-C479|Peripheral_Nerve|880|Sarcoma|8800/3|Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C470-C476,C478-C479|Peripheral_Nerve|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C470-C476,C478-C479|Peripheral_Nerve|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C470-C476,C478-C479|Peripheral_Nerve|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C470-C476,C478-C479|Peripheral_Nerve|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C470-C476,C478-C479|Peripheral_Nerve|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C470-C476,C478-C479|Peripheral_Nerve|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C470-C476,C478-C479|Peripheral_Nerve|882|Sarcoma|8825/3|Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C470-C476,C478-C479|Peripheral_Nerve|883|Benign_Fibrous_Histiocytoma|8832/3|Dermatofibrosarcoma_Protuberans
C470-C476,C478-C479|Peripheral_Nerve|883|Benign_Fibrous_Histiocytoma|8833/3|Dermatofibrosarcoma_Protuberans
C470-C476,C478-C479|Peripheral_Nerve|884|Myxosarcoma|8840/3|Myxosarcoma
C470-C476,C478-C479|Peripheral_Nerve|885|Liposarcoma|8850/3|Liposarcoma
C470-C476,C478-C479|Peripheral_Nerve|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C470-C476,C478-C479|Peripheral_Nerve|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C470-C476,C478-C479|Peripheral_Nerve|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C470-C476,C478-C479|Peripheral_Nerve|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C470-C476,C478-C479|Peripheral_Nerve|885|Liposarcoma|8855/3|Liposarcoma
C470-C476,C478-C479|Peripheral_Nerve|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C470-C476,C478-C479|Peripheral_Nerve|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C470-C476,C478-C479|Peripheral_Nerve|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C470-C476,C478-C479|Peripheral_Nerve|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C470-C476,C478-C479|Peripheral_Nerve|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C470-C476,C478-C479|Peripheral_Nerve|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C470-C476,C478-C479|Peripheral_Nerve|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C470-C476,C478-C479|Peripheral_Nerve|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|904|Synovial_Sarcoma|9040/3|Synovial_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|904|Synovial_Sarcoma|9041/3|Spindle_Cell_Synovial_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|904|Synovial_Sarcoma|9042/3|Epithelial_Synovial_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|904|Synovial_Sarcoma|9043/3|Biphasic_Synovial_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|904|Synovial_Sarcoma|9044/3|Clear_Cell_Sarcoma_Of_Soft_Tissue_C0206651
C470-C476,C478-C479|Peripheral_Nerve|908|Teratoma|9080/3|Immature_Teratoma
C470-C476,C478-C479|Peripheral_Nerve|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C470-C476,C478-C479|Peripheral_Nerve|908|Teratoma|9082/3|Immature_Teratoma
C470-C476,C478-C479|Peripheral_Nerve|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C470-C476,C478-C479|Peripheral_Nerve|908|Teratoma|9084/3|Teratoma
C470-C476,C478-C479|Peripheral_Nerve|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C470-C476,C478-C479|Peripheral_Nerve|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C470-C476,C478-C479|Peripheral_Nerve|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C470-C476,C478-C479|Peripheral_Nerve|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C470-C476,C478-C479|Peripheral_Nerve|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C470-C476,C478-C479|Peripheral_Nerve|917|Lymphangiosarcoma|9170/3|Lymphangiosarcoma
C470-C476,C478-C479|Peripheral_Nerve|924|Neoplasm|9240/3|Mesenchymal_Chondrosarcoma
C470-C476,C478-C479|Peripheral_Nerve|924|Neoplasm|9242/3|Clear_Cell_Chondrosarcoma
C470-C476,C478-C479|Peripheral_Nerve|924|Neoplasm|9243/3|Dedifferentiated_Chondrosarcoma
C470-C476,C478-C479|Peripheral_Nerve|925|Bone_Neoplasm|9251/3|Giant_Cell_Tumor_Of_Soft_Tissue
C470-C476,C478-C479|Peripheral_Nerve|925|Bone_Neoplasm|9252/3|Malignant_Tenosynovial_Giant_Cell_Tumor
C470-C476,C478-C479|Peripheral_Nerve|936|Neuroepithelioma__Peripheral|9364/3|Neuroepithelioma__Peripheral
C470-C476,C478-C479|Peripheral_Nerve|936|Neuroepithelioma__Peripheral|9365/3|Askin_Tumor
C470-C476,C478-C479|Peripheral_Nerve|937|Chordoma|9370/3|Chordoma
C470-C476,C478-C479|Peripheral_Nerve|937|Chordoma|9371/3|Chondroid_Chordoma
C470-C476,C478-C479|Peripheral_Nerve|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C470-C476,C478-C479|Peripheral_Nerve|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C470-C476,C478-C479|Peripheral_Nerve|950|Neuroblastoma|9500/3|Neuroblastoma
C470-C476,C478-C479|Peripheral_Nerve|950|Neuroblastoma|9501/3|Medulloepithelioma
C470-C476,C478-C479|Peripheral_Nerve|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C470-C476,C478-C479|Peripheral_Nerve|950|Neuroblastoma|9503/3|Neuroepithelioma
C470-C476,C478-C479|Peripheral_Nerve|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C470-C476,C478-C479|Peripheral_Nerve|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C470-C476,C478-C479|Peripheral_Nerve|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C470-C476,C478-C479|Peripheral_Nerve|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9542/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C470-C476,C478-C479|Peripheral_Nerve|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C470-C476,C478-C479|Peripheral_Nerve|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C470-C476,C478-C479|Peripheral_Nerve|957|Perineurioma|9571/3|Malignant_Perineurioma
C470-C476,C478-C479|Peripheral_Nerve|958|Granular_Cell_Tumor|9580/3|Malignant_Granular_Cell_Tumor
C470-C476,C478-C479|Peripheral_Nerve|958|Granular_Cell_Tumor|9581/3|Alveolar_Soft_Part_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|959|Lymphoma|9590/3|Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C470-C476,C478-C479|Peripheral_Nerve|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C470-C476,C478-C479|Peripheral_Nerve|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C470-C476,C478-C479|Peripheral_Nerve|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C470-C476,C478-C479|Peripheral_Nerve|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C470-C476,C478-C479|Peripheral_Nerve|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C470-C476,C478-C479|Peripheral_Nerve|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C470-C476,C478-C479|Peripheral_Nerve|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C470-C476,C478-C479|Peripheral_Nerve|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C470-C476,C478-C479|Peripheral_Nerve|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C470-C476,C478-C479|Peripheral_Nerve|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C470-C476,C478-C479|Peripheral_Nerve|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C470-C476,C478-C479|Peripheral_Nerve|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C470-C476,C478-C479|Peripheral_Nerve|972|Lymphoblastic_Lymphoma|9726/3|T_Cell_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|973|Plasmacytoma|9731/3|Plasmacytoma
C470-C476,C478-C479|Peripheral_Nerve|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C470-C476,C478-C479|Peripheral_Nerve|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C470-C476,C478-C479|Peripheral_Nerve|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C470-C476,C478-C479|Peripheral_Nerve|975|Neoplasm|9750/3|Malignant_Histiocytosis
C470-C476,C478-C479|Peripheral_Nerve|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C470-C476,C478-C479|Peripheral_Nerve|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C470-C476,C478-C479|Peripheral_Nerve|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C470-C476,C478-C479|Peripheral_Nerve|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9812/3|Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9813/3|Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9814/3|Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9816/3|Hypodiploid_ALL
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9817/3|Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9818/3|Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|981|Neoplasm|9819/3|Leukemia__B_Cell
C470-C476,C478-C479|Peripheral_Nerve|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C470-C476,C478-C479|Peripheral_Nerve|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C470-C476,C478-C479|Peripheral_Nerve|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C470-C476,C478-C479|Peripheral_Nerve|993|Myeloid_Sarcoma|9930/3|Myeloid_Sarcoma
C470-C476,C478-C479|Peripheral_Nerve|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C470-C476,C478-C479|Peripheral_Nerve|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C470-C476,C478-C479|Peripheral_Nerve|997|Neoplasm|9971/3|Polymorphic_PTLD
C470-C476,C478-C479|Peripheral_Nerve|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C480-C482,C488|Retroperitoneal_Space|800|Neoplasm|8000/3|Malignant_Neoplasm
C480-C482,C488|Retroperitoneal_Space|800|Neoplasm|8001/3|Malignant_Cell
C480-C482,C488|Retroperitoneal_Space|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C480-C482,C488|Retroperitoneal_Space|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C480-C482,C488|Retroperitoneal_Space|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C480-C482,C488|Retroperitoneal_Space|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C480-C482,C488|Retroperitoneal_Space|846|Papillary_Serous_Cystadenocarcinoma|8461/3|Serous_Surface_Papillary_Carcinoma
C480-C482,C488|Retroperitoneal_Space|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C480-C482,C488|Retroperitoneal_Space|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C480-C482,C488|Retroperitoneal_Space|871|Malignant_Glomus_Tumor|8714/3|Malignant_PEComa
C480-C482,C488|Retroperitoneal_Space|880|Sarcoma|8800/3|Sarcoma
C480-C482,C488|Retroperitoneal_Space|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C480-C482,C488|Retroperitoneal_Space|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C480-C482,C488|Retroperitoneal_Space|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C480-C482,C488|Retroperitoneal_Space|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C480-C482,C488|Retroperitoneal_Space|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C480-C482,C488|Retroperitoneal_Space|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C480-C482,C488|Retroperitoneal_Space|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C480-C482,C488|Retroperitoneal_Space|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C480-C482,C488|Retroperitoneal_Space|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C480-C482,C488|Retroperitoneal_Space|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C480-C482,C488|Retroperitoneal_Space|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C480-C482,C488|Retroperitoneal_Space|882|Sarcoma|8825/3|Sarcoma
C480-C482,C488|Retroperitoneal_Space|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C480-C482,C488|Retroperitoneal_Space|884|Myxosarcoma|8840/3|Myxosarcoma
C480-C482,C488|Retroperitoneal_Space|885|Liposarcoma|8850/3|Liposarcoma
C480-C482,C488|Retroperitoneal_Space|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C480-C482,C488|Retroperitoneal_Space|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C480-C482,C488|Retroperitoneal_Space|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C480-C482,C488|Retroperitoneal_Space|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C480-C482,C488|Retroperitoneal_Space|885|Liposarcoma|8855/3|Liposarcoma
C480-C482,C488|Retroperitoneal_Space|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C480-C482,C488|Retroperitoneal_Space|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C480-C482,C488|Retroperitoneal_Space|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C480-C482,C488|Retroperitoneal_Space|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C480-C482,C488|Retroperitoneal_Space|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C480-C482,C488|Retroperitoneal_Space|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C480-C482,C488|Retroperitoneal_Space|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C480-C482,C488|Retroperitoneal_Space|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C480-C482,C488|Retroperitoneal_Space|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C480-C482,C488|Retroperitoneal_Space|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C480-C482,C488|Retroperitoneal_Space|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C480-C482,C488|Retroperitoneal_Space|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C480-C482,C488|Retroperitoneal_Space|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C480-C482,C488|Retroperitoneal_Space|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C480-C482,C488|Retroperitoneal_Space|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C480-C482,C488|Retroperitoneal_Space|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C480-C482,C488|Retroperitoneal_Space|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C480-C482,C488|Retroperitoneal_Space|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C480-C482,C488|Retroperitoneal_Space|905|Malignant_Mesothelioma|9050/3|Malignant_Mesothelioma
C480-C482,C488|Retroperitoneal_Space|905|Malignant_Mesothelioma|9051/3|Sarcomatoid_Mesothelioma
C480-C482,C488|Retroperitoneal_Space|905|Malignant_Mesothelioma|9052/3|Mesothelioma
C480-C482,C488|Retroperitoneal_Space|905|Malignant_Mesothelioma|9053/3|Biphasic_Mesothelioma
C480-C482,C488|Retroperitoneal_Space|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C480-C482,C488|Retroperitoneal_Space|906|Germ_Cell_Tumor|9064/3|Germinoma
C480-C482,C488|Retroperitoneal_Space|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C480-C482,C488|Retroperitoneal_Space|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C480-C482,C488|Retroperitoneal_Space|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C480-C482,C488|Retroperitoneal_Space|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C480-C482,C488|Retroperitoneal_Space|908|Teratoma|9080/3|Immature_Teratoma
C480-C482,C488|Retroperitoneal_Space|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C480-C482,C488|Retroperitoneal_Space|908|Teratoma|9082/3|Immature_Teratoma
C480-C482,C488|Retroperitoneal_Space|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C480-C482,C488|Retroperitoneal_Space|908|Teratoma|9084/3|Teratoma
C480-C482,C488|Retroperitoneal_Space|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C480-C482,C488|Retroperitoneal_Space|911|Mesonephroma|9110/3|Mesonephroma
C480-C482,C488|Retroperitoneal_Space|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C480-C482,C488|Retroperitoneal_Space|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C480-C482,C488|Retroperitoneal_Space|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C480-C482,C488|Retroperitoneal_Space|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C480-C482,C488|Retroperitoneal_Space|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C480-C482,C488|Retroperitoneal_Space|950|Neuroblastoma|9500/3|Neuroblastoma
C480-C482,C488|Retroperitoneal_Space|950|Neuroblastoma|9501/3|Medulloepithelioma
C480-C482,C488|Retroperitoneal_Space|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C480-C482,C488|Retroperitoneal_Space|950|Neuroblastoma|9503/3|Neuroepithelioma
C480-C482,C488|Retroperitoneal_Space|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C480-C482,C488|Retroperitoneal_Space|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C480-C482,C488|Retroperitoneal_Space|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C480-C482,C488|Retroperitoneal_Space|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C480-C482,C488|Retroperitoneal_Space|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C480-C482,C488|Retroperitoneal_Space|957|Perineurioma|9571/3|Malignant_Perineurioma
C480-C482,C488|Retroperitoneal_Space|959|Lymphoma|9590/3|Lymphoma
C480-C482,C488|Retroperitoneal_Space|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C480-C482,C488|Retroperitoneal_Space|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C480-C482,C488|Retroperitoneal_Space|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C480-C482,C488|Retroperitoneal_Space|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C480-C482,C488|Retroperitoneal_Space|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C480-C482,C488|Retroperitoneal_Space|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C480-C482,C488|Retroperitoneal_Space|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C480-C482,C488|Retroperitoneal_Space|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C480-C482,C488|Retroperitoneal_Space|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C480-C482,C488|Retroperitoneal_Space|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C480-C482,C488|Retroperitoneal_Space|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C480-C482,C488|Retroperitoneal_Space|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C480-C482,C488|Retroperitoneal_Space|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C480-C482,C488|Retroperitoneal_Space|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C480-C482,C488|Retroperitoneal_Space|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C480-C482,C488|Retroperitoneal_Space|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C480-C482,C488|Retroperitoneal_Space|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C480-C482,C488|Retroperitoneal_Space|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C480-C482,C488|Retroperitoneal_Space|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C480-C482,C488|Retroperitoneal_Space|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C480-C482,C488|Retroperitoneal_Space|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C480-C482,C488|Retroperitoneal_Space|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C480-C482,C488|Retroperitoneal_Space|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C480-C482,C488|Retroperitoneal_Space|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C480-C482,C488|Retroperitoneal_Space|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C480-C482,C488|Retroperitoneal_Space|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C480-C482,C488|Retroperitoneal_Space|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C480-C482,C488|Retroperitoneal_Space|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C480-C482,C488|Retroperitoneal_Space|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C480-C482,C488|Retroperitoneal_Space|973|Plasmacytoma|9731/3|Plasmacytoma
C480-C482,C488|Retroperitoneal_Space|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C480-C482,C488|Retroperitoneal_Space|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C480-C482,C488|Retroperitoneal_Space|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C480-C482,C488|Retroperitoneal_Space|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C480-C482,C488|Retroperitoneal_Space|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C480-C482,C488|Retroperitoneal_Space|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C480-C482,C488|Retroperitoneal_Space|975|Neoplasm|9750/3|Malignant_Histiocytosis
C480-C482,C488|Retroperitoneal_Space|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C480-C482,C488|Retroperitoneal_Space|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C480-C482,C488|Retroperitoneal_Space|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C480-C482,C488|Retroperitoneal_Space|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C480-C482,C488|Retroperitoneal_Space|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C480-C482,C488|Retroperitoneal_Space|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C480-C482,C488|Retroperitoneal_Space|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C480-C482,C488|Retroperitoneal_Space|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9812/3|Lymphoma
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9813/3|Lymphoma
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9814/3|Lymphoma
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9816/3|Hypodiploid_ALL
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9817/3|Lymphoma
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9818/3|Lymphoma
C480-C482,C488|Retroperitoneal_Space|981|Neoplasm|9819/3|Leukemia__B_Cell
C480-C482,C488|Retroperitoneal_Space|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C480-C482,C488|Retroperitoneal_Space|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C480-C482,C488|Retroperitoneal_Space|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C480-C482,C488|Retroperitoneal_Space|993|Myeloid_Sarcoma|9930/3|Myeloid_Sarcoma
C480-C482,C488|Retroperitoneal_Space|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C480-C482,C488|Retroperitoneal_Space|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C480-C482,C488|Retroperitoneal_Space|997|Neoplasm|9971/3|Polymorphic_PTLD
C480-C482,C488|Retroperitoneal_Space|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C490-C496,C498-C499|Body_Tissue|800|Neoplasm|8000/3|Malignant_Neoplasm
C490-C496,C498-C499|Body_Tissue|800|Neoplasm|8001/3|Malignant_Cell
C490-C496,C498-C499|Body_Tissue|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C490-C496,C498-C499|Body_Tissue|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C490-C496,C498-C499|Body_Tissue|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C490-C496,C498-C499|Body_Tissue|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C490-C496,C498-C499|Body_Tissue|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C490-C496,C498-C499|Body_Tissue|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C490-C496,C498-C499|Body_Tissue|880|Sarcoma|8800/3|Sarcoma
C490-C496,C498-C499|Body_Tissue|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C490-C496,C498-C499|Body_Tissue|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C490-C496,C498-C499|Body_Tissue|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C490-C496,C498-C499|Body_Tissue|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C490-C496,C498-C499|Body_Tissue|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C490-C496,C498-C499|Body_Tissue|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C490-C496,C498-C499|Body_Tissue|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C490-C496,C498-C499|Body_Tissue|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C490-C496,C498-C499|Body_Tissue|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C490-C496,C498-C499|Body_Tissue|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C490-C496,C498-C499|Body_Tissue|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C490-C496,C498-C499|Body_Tissue|882|Sarcoma|8825/3|Sarcoma
C490-C496,C498-C499|Body_Tissue|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C490-C496,C498-C499|Body_Tissue|883|Benign_Fibrous_Histiocytoma|8832/3|Dermatofibrosarcoma_Protuberans
C490-C496,C498-C499|Body_Tissue|883|Benign_Fibrous_Histiocytoma|8833/3|Dermatofibrosarcoma_Protuberans
C490-C496,C498-C499|Body_Tissue|884|Myxosarcoma|8840/3|Myxosarcoma
C490-C496,C498-C499|Body_Tissue|884|Myxosarcoma|8842/3|Sarcoma
C490-C496,C498-C499|Body_Tissue|885|Liposarcoma|8850/3|Liposarcoma
C490-C496,C498-C499|Body_Tissue|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C490-C496,C498-C499|Body_Tissue|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C490-C496,C498-C499|Body_Tissue|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C490-C496,C498-C499|Body_Tissue|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C490-C496,C498-C499|Body_Tissue|885|Liposarcoma|8855/3|Liposarcoma
C490-C496,C498-C499|Body_Tissue|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C490-C496,C498-C499|Body_Tissue|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C490-C496,C498-C499|Body_Tissue|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C490-C496,C498-C499|Body_Tissue|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C490-C496,C498-C499|Body_Tissue|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C490-C496,C498-C499|Body_Tissue|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C490-C496,C498-C499|Body_Tissue|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C490-C496,C498-C499|Body_Tissue|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C490-C496,C498-C499|Body_Tissue|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C490-C496,C498-C499|Body_Tissue|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C490-C496,C498-C499|Body_Tissue|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C490-C496,C498-C499|Body_Tissue|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C490-C496,C498-C499|Body_Tissue|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C490-C496,C498-C499|Body_Tissue|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C490-C496,C498-C499|Body_Tissue|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C490-C496,C498-C499|Body_Tissue|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C490-C496,C498-C499|Body_Tissue|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C490-C496,C498-C499|Body_Tissue|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C490-C496,C498-C499|Body_Tissue|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C490-C496,C498-C499|Body_Tissue|904|Synovial_Sarcoma|9040/3|Synovial_Sarcoma
C490-C496,C498-C499|Body_Tissue|904|Synovial_Sarcoma|9041/3|Spindle_Cell_Synovial_Sarcoma
C490-C496,C498-C499|Body_Tissue|904|Synovial_Sarcoma|9042/3|Epithelial_Synovial_Sarcoma
C490-C496,C498-C499|Body_Tissue|904|Synovial_Sarcoma|9043/3|Biphasic_Synovial_Sarcoma
C490-C496,C498-C499|Body_Tissue|904|Synovial_Sarcoma|9044/3|Clear_Cell_Sarcoma_Of_Soft_Tissue_C0206651
C490-C496,C498-C499|Body_Tissue|908|Teratoma|9080/3|Immature_Teratoma
C490-C496,C498-C499|Body_Tissue|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C490-C496,C498-C499|Body_Tissue|908|Teratoma|9082/3|Immature_Teratoma
C490-C496,C498-C499|Body_Tissue|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C490-C496,C498-C499|Body_Tissue|908|Teratoma|9084/3|Teratoma
C490-C496,C498-C499|Body_Tissue|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C490-C496,C498-C499|Body_Tissue|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C490-C496,C498-C499|Body_Tissue|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C490-C496,C498-C499|Body_Tissue|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C490-C496,C498-C499|Body_Tissue|913|Hemangioendothelioma|9137/3|Intimal_Sarcoma
C490-C496,C498-C499|Body_Tissue|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C490-C496,C498-C499|Body_Tissue|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C490-C496,C498-C499|Body_Tissue|917|Lymphangiosarcoma|9170/3|Lymphangiosarcoma
C490-C496,C498-C499|Body_Tissue|924|Neoplasm|9240/3|Mesenchymal_Chondrosarcoma
C490-C496,C498-C499|Body_Tissue|924|Neoplasm|9242/3|Clear_Cell_Chondrosarcoma
C490-C496,C498-C499|Body_Tissue|924|Neoplasm|9243/3|Dedifferentiated_Chondrosarcoma
C490-C496,C498-C499|Body_Tissue|925|Bone_Neoplasm|9251/3|Giant_Cell_Tumor_Of_Soft_Tissue
C490-C496,C498-C499|Body_Tissue|925|Bone_Neoplasm|9252/3|Malignant_Tenosynovial_Giant_Cell_Tumor
C490-C496,C498-C499|Body_Tissue|936|Neuroepithelioma__Peripheral|9364/3|Neuroepithelioma__Peripheral
C490-C496,C498-C499|Body_Tissue|936|Neuroepithelioma__Peripheral|9365/3|Askin_Tumor
C490-C496,C498-C499|Body_Tissue|937|Chordoma|9370/3|Chordoma
C490-C496,C498-C499|Body_Tissue|937|Chordoma|9371/3|Chondroid_Chordoma
C490-C496,C498-C499|Body_Tissue|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C490-C496,C498-C499|Body_Tissue|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C490-C496,C498-C499|Body_Tissue|950|Neuroblastoma|9500/3|Neuroblastoma
C490-C496,C498-C499|Body_Tissue|950|Neuroblastoma|9501/3|Medulloepithelioma
C490-C496,C498-C499|Body_Tissue|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C490-C496,C498-C499|Body_Tissue|950|Neuroblastoma|9503/3|Neuroepithelioma
C490-C496,C498-C499|Body_Tissue|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C490-C496,C498-C499|Body_Tissue|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C490-C496,C498-C499|Body_Tissue|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C490-C496,C498-C499|Body_Tissue|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C490-C496,C498-C499|Body_Tissue|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C490-C496,C498-C499|Body_Tissue|957|Perineurioma|9571/3|Malignant_Perineurioma
C490-C496,C498-C499|Body_Tissue|958|Granular_Cell_Tumor|9580/3|Malignant_Granular_Cell_Tumor
C490-C496,C498-C499|Body_Tissue|958|Granular_Cell_Tumor|9581/3|Alveolar_Soft_Part_Sarcoma
C490-C496,C498-C499|Body_Tissue|959|Lymphoma|9590/3|Lymphoma
C490-C496,C498-C499|Body_Tissue|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C490-C496,C498-C499|Body_Tissue|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C490-C496,C498-C499|Body_Tissue|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C490-C496,C498-C499|Body_Tissue|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C490-C496,C498-C499|Body_Tissue|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C490-C496,C498-C499|Body_Tissue|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C490-C496,C498-C499|Body_Tissue|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C490-C496,C498-C499|Body_Tissue|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C490-C496,C498-C499|Body_Tissue|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C490-C496,C498-C499|Body_Tissue|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C490-C496,C498-C499|Body_Tissue|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C490-C496,C498-C499|Body_Tissue|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C490-C496,C498-C499|Body_Tissue|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C490-C496,C498-C499|Body_Tissue|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C490-C496,C498-C499|Body_Tissue|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C490-C496,C498-C499|Body_Tissue|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C490-C496,C498-C499|Body_Tissue|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C490-C496,C498-C499|Body_Tissue|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C490-C496,C498-C499|Body_Tissue|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C490-C496,C498-C499|Body_Tissue|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C490-C496,C498-C499|Body_Tissue|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C490-C496,C498-C499|Body_Tissue|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C490-C496,C498-C499|Body_Tissue|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C490-C496,C498-C499|Body_Tissue|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C490-C496,C498-C499|Body_Tissue|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C490-C496,C498-C499|Body_Tissue|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C490-C496,C498-C499|Body_Tissue|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C490-C496,C498-C499|Body_Tissue|972|Lymphoblastic_Lymphoma|9726/3|T_Cell_Lymphoma
C490-C496,C498-C499|Body_Tissue|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C490-C496,C498-C499|Body_Tissue|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C490-C496,C498-C499|Body_Tissue|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C490-C496,C498-C499|Body_Tissue|973|Plasmacytoma|9731/3|Plasmacytoma
C490-C496,C498-C499|Body_Tissue|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C490-C496,C498-C499|Body_Tissue|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C490-C496,C498-C499|Body_Tissue|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C490-C496,C498-C499|Body_Tissue|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C490-C496,C498-C499|Body_Tissue|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C490-C496,C498-C499|Body_Tissue|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C490-C496,C498-C499|Body_Tissue|975|Neoplasm|9750/3|Malignant_Histiocytosis
C490-C496,C498-C499|Body_Tissue|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C490-C496,C498-C499|Body_Tissue|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C490-C496,C498-C499|Body_Tissue|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C490-C496,C498-C499|Body_Tissue|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C490-C496,C498-C499|Body_Tissue|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C490-C496,C498-C499|Body_Tissue|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C490-C496,C498-C499|Body_Tissue|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C490-C496,C498-C499|Body_Tissue|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9812/3|Lymphoma
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9813/3|Lymphoma
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9814/3|Lymphoma
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9816/3|Hypodiploid_ALL
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9817/3|Lymphoma
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9818/3|Lymphoma
C490-C496,C498-C499|Body_Tissue|981|Neoplasm|9819/3|Leukemia__B_Cell
C490-C496,C498-C499|Body_Tissue|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C490-C496,C498-C499|Body_Tissue|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C490-C496,C498-C499|Body_Tissue|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C490-C496,C498-C499|Body_Tissue|993|Myeloid_Sarcoma|9930/3|Myeloid_Sarcoma
C490-C496,C498-C499|Body_Tissue|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C490-C496,C498-C499|Body_Tissue|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C490-C496,C498-C499|Body_Tissue|997|Neoplasm|9971/3|Polymorphic_PTLD
C490-C496,C498-C499|Body_Tissue|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C500-C506,C508-C509|Breast|800|Neoplasm|8000/3|Malignant_Neoplasm
C500-C506,C508-C509|Breast|800|Neoplasm|8001/3|Malignant_Cell
C500-C506,C508-C509|Breast|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C500-C506,C508-C509|Breast|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C500-C506,C508-C509|Breast|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C500-C506,C508-C509|Breast|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C500-C506,C508-C509|Breast|801|Carcinoma|8010/2|In_Situ_Cancer
C500-C506,C508-C509|Breast|801|Carcinoma|8010/3|Carcinoma
C500-C506,C508-C509|Breast|801|Carcinoma|8011/3|Malignant_Epithelioma
C500-C506,C508-C509|Breast|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C500-C506,C508-C509|Breast|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C500-C506,C508-C509|Breast|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C500-C506,C508-C509|Breast|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C500-C506,C508-C509|Breast|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C500-C506,C508-C509|Breast|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C500-C506,C508-C509|Breast|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C500-C506,C508-C509|Breast|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C500-C506,C508-C509|Breast|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C500-C506,C508-C509|Breast|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C500-C506,C508-C509|Breast|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C500-C506,C508-C509|Breast|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C500-C506,C508-C509|Breast|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C500-C506,C508-C509|Breast|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C500-C506,C508-C509|Breast|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C500-C506,C508-C509|Breast|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C500-C506,C508-C509|Breast|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C500-C506,C508-C509|Breast|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C500-C506,C508-C509|Breast|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C500-C506,C508-C509|Breast|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C500-C506,C508-C509|Breast|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8140/3|Adenocarcinoma
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C500-C506,C508-C509|Breast|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C500-C506,C508-C509|Breast|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C500-C506,C508-C509|Breast|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C500-C506,C508-C509|Breast|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C500-C506,C508-C509|Breast|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C500-C506,C508-C509|Breast|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C500-C506,C508-C509|Breast|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C500-C506,C508-C509|Breast|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C500-C506,C508-C509|Breast|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C500-C506,C508-C509|Breast|825|Bronchioloalveolar_Adenocarcinoma|8251/3|Bronchioloalveolar_Adenocarcinoma
C500-C506,C508-C509|Breast|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C500-C506,C508-C509|Breast|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C500-C506,C508-C509|Breast|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C500-C506,C508-C509|Breast|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C500-C506,C508-C509|Breast|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C500-C506,C508-C509|Breast|831|Clear_Cell_Adenocarcinoma|8314/3|Lipid_Rich_Carcinoma
C500-C506,C508-C509|Breast|831|Clear_Cell_Adenocarcinoma|8315/3|Glycogen_Rich_Carcinoma
C500-C506,C508-C509|Breast|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C500-C506,C508-C509|Breast|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C500-C506,C508-C509|Breast|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C500-C506,C508-C509|Breast|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C500-C506,C508-C509|Breast|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C500-C506,C508-C509|Breast|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C500-C506,C508-C509|Breast|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8500/1|Ductal_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8500/2|Ductal_Breast_Carcinoma_In_Situ
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8500/3|Invasive_Breast_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8501/2|Comedocarcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8501/3|Comedocarcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8502/3|Secretory_Breast_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8503/2|Intraductal_Papillary_Breast_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8503/3|Intraductal_Papillary_Breast_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8504/2|Intracystic_Papillary_Breast_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8504/3|Intracystic_Papillary_Breast_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8507/2|Micropapillary_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8507/3|Micropapillary_Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8508/3|Carcinoma
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8509/2|Solid_Papillary_Carcinoma_In_Situ
C500-C506,C508-C509|Breast|850|Ductal_Carcinoma|8509/3|Papillary_Carcinoma
C500-C506,C508-C509|Breast|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C500-C506,C508-C509|Breast|851|Medullary_Carcinoma|8512/3|Medullary_Carcinoma
C500-C506,C508-C509|Breast|851|Medullary_Carcinoma|8513/3|Medullary_Carcinoma
C500-C506,C508-C509|Breast|851|Medullary_Carcinoma|8514/3|Ductal_Carcinoma
C500-C506,C508-C509|Breast|851|Medullary_Carcinoma|8519/2|Pleomorphic_Lobular_Carcinoma_In_Situ
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8520/2|Lobular_Breast_Carcinoma_In_Situ
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8520/3|Carcinoma__Lobular
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8521/3|Invasive_Ductal_Breast_Carcinoma
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8522/2|Carcinoma
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8522/3|Intraductal_And_Lobular_Carcinoma
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8523/2|Carcinoma
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8523/3|Carcinoma
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8524/3|Invasive_Lobular_Breast_Carcinoma
C500-C506,C508-C509|Breast|852|Intraductal_And_Lobular_Carcinoma|8525/3|Terminal_Duct_Adenocarcinoma
C500-C506,C508-C509|Breast|853|Inflammatory_Carcinoma|8530/3|Inflammatory_Carcinoma
C500-C506,C508-C509|Breast|854|Paget_s_Disease__Mammary|8540/3|Paget_s_Disease__Mammary
C500-C506,C508-C509|Breast|854|Paget_s_Disease__Mammary|8541/3|Ductal_Carcinoma
C500-C506,C508-C509|Breast|854|Paget_s_Disease__Mammary|8543/3|Paget_Disease
C500-C506,C508-C509|Breast|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C500-C506,C508-C509|Breast|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C500-C506,C508-C509|Breast|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C500-C506,C508-C509|Breast|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C500-C506,C508-C509|Breast|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C500-C506,C508-C509|Breast|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C500-C506,C508-C509|Breast|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C500-C506,C508-C509|Breast|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C500-C506,C508-C509|Breast|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C500-C506,C508-C509|Breast|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C500-C506,C508-C509|Breast|880|Sarcoma|8800/3|Sarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C500-C506,C508-C509|Breast|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C500-C506,C508-C509|Breast|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C500-C506,C508-C509|Breast|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C500-C506,C508-C509|Breast|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C500-C506,C508-C509|Breast|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C500-C506,C508-C509|Breast|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C500-C506,C508-C509|Breast|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C500-C506,C508-C509|Breast|882|Sarcoma|8825/3|Sarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8850/3|Liposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C500-C506,C508-C509|Breast|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8855/3|Liposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C500-C506,C508-C509|Breast|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C500-C506,C508-C509|Breast|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C500-C506,C508-C509|Breast|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C500-C506,C508-C509|Breast|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C500-C506,C508-C509|Breast|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C500-C506,C508-C509|Breast|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C500-C506,C508-C509|Breast|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C500-C506,C508-C509|Breast|898|Carcinosarcoma|8980/3|Carcinosarcoma
C500-C506,C508-C509|Breast|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C500-C506,C508-C509|Breast|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C500-C506,C508-C509|Breast|898|Carcinosarcoma|8983/3|Adenomyoepithelioma_With_Carcinoma
C500-C506,C508-C509|Breast|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C500-C506,C508-C509|Breast|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C500-C506,C508-C509|Breast|902|Phyllodes_Tumor|9020/3|Malignant_Phyllodes_Tumor
C500-C506,C508-C509|Breast|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C500-C506,C508-C509|Breast|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C500-C506,C508-C509|Breast|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C500-C506,C508-C509|Breast|958|Granular_Cell_Tumor|9580/3|Malignant_Granular_Cell_Tumor
C500-C506,C508-C509|Breast|958|Granular_Cell_Tumor|9581/3|Alveolar_Soft_Part_Sarcoma
C500-C506,C508-C509|Breast|959|Lymphoma|9590/3|Lymphoma
C500-C506,C508-C509|Breast|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C500-C506,C508-C509|Breast|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C500-C506,C508-C509|Breast|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C500-C506,C508-C509|Breast|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C500-C506,C508-C509|Breast|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C500-C506,C508-C509|Breast|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C500-C506,C508-C509|Breast|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C500-C506,C508-C509|Breast|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C500-C506,C508-C509|Breast|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C500-C506,C508-C509|Breast|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C500-C506,C508-C509|Breast|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C500-C506,C508-C509|Breast|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C500-C506,C508-C509|Breast|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C500-C506,C508-C509|Breast|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C500-C506,C508-C509|Breast|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C500-C506,C508-C509|Breast|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C500-C506,C508-C509|Breast|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C500-C506,C508-C509|Breast|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C500-C506,C508-C509|Breast|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C500-C506,C508-C509|Breast|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C500-C506,C508-C509|Breast|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C500-C506,C508-C509|Breast|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C500-C506,C508-C509|Breast|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C500-C506,C508-C509|Breast|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C500-C506,C508-C509|Breast|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C500-C506,C508-C509|Breast|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C500-C506,C508-C509|Breast|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C500-C506,C508-C509|Breast|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C500-C506,C508-C509|Breast|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9731/3|Plasmacytoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C500-C506,C508-C509|Breast|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C500-C506,C508-C509|Breast|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C500-C506,C508-C509|Breast|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C500-C506,C508-C509|Breast|975|Neoplasm|9750/3|Malignant_Histiocytosis
C500-C506,C508-C509|Breast|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C500-C506,C508-C509|Breast|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C500-C506,C508-C509|Breast|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C500-C506,C508-C509|Breast|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C500-C506,C508-C509|Breast|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C500-C506,C508-C509|Breast|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C500-C506,C508-C509|Breast|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C500-C506,C508-C509|Breast|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C500-C506,C508-C509|Breast|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C500-C506,C508-C509|Breast|981|Neoplasm|9812/3|Lymphoma
C500-C506,C508-C509|Breast|981|Neoplasm|9813/3|Lymphoma
C500-C506,C508-C509|Breast|981|Neoplasm|9814/3|Lymphoma
C500-C506,C508-C509|Breast|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C500-C506,C508-C509|Breast|981|Neoplasm|9816/3|Hypodiploid_ALL
C500-C506,C508-C509|Breast|981|Neoplasm|9817/3|Lymphoma
C500-C506,C508-C509|Breast|981|Neoplasm|9818/3|Lymphoma
C500-C506,C508-C509|Breast|981|Neoplasm|9819/3|Leukemia__B_Cell
C500-C506,C508-C509|Breast|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C500-C506,C508-C509|Breast|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C500-C506,C508-C509|Breast|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C500-C506,C508-C509|Breast|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C500-C506,C508-C509|Breast|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C500-C506,C508-C509|Breast|997|Neoplasm|9971/3|Polymorphic_PTLD
C500-C506,C508-C509|Breast|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C510-C512,C518, C529|Vagina|800|Neoplasm|8000/3|Malignant_Neoplasm
C510-C512,C518, C529|Vagina|800|Neoplasm|8001/3|Malignant_Cell
C510-C512,C518, C529|Vagina|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C510-C512,C518, C529|Vagina|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C510-C512,C518, C529|Vagina|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C510-C512,C518, C529|Vagina|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C510-C512,C518, C529|Vagina|801|Carcinoma|8010/2|In_Situ_Cancer
C510-C512,C518, C529|Vagina|801|Carcinoma|8010/3|Carcinoma
C510-C512,C518, C529|Vagina|801|Carcinoma|8011/3|Malignant_Epithelioma
C510-C512,C518, C529|Vagina|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C510-C512,C518, C529|Vagina|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C510-C512,C518, C529|Vagina|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C510-C512,C518, C529|Vagina|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C510-C512,C518, C529|Vagina|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C510-C512,C518, C529|Vagina|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C510-C512,C518, C529|Vagina|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C510-C512,C518, C529|Vagina|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C510-C512,C518, C529|Vagina|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C510-C512,C518, C529|Vagina|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C510-C512,C518, C529|Vagina|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8071/2|Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8077/2|Intraepithelial_Neoplasia
C510-C512,C518, C529|Vagina|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C510-C512,C518, C529|Vagina|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C510-C512,C518, C529|Vagina|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|809|Basal_Cell_Carcinoma|8090/3|Basal_Cell_Carcinoma
C510-C512,C518, C529|Vagina|809|Basal_Cell_Carcinoma|8091/3|Superficial_Basal_Cell_Carcinoma
C510-C512,C518, C529|Vagina|809|Basal_Cell_Carcinoma|8092/3|Skin_Infiltrating_Basal_Cell_Carcinoma
C510-C512,C518, C529|Vagina|809|Basal_Cell_Carcinoma|8093/3|Fibroepithelioma_Of_Pinkus
C510-C512,C518, C529|Vagina|809|Basal_Cell_Carcinoma|8094/3|Skin_Basosquamous_Cell_Carcinoma
C510-C512,C518, C529|Vagina|809|Basal_Cell_Carcinoma|8095/3|Skin_Metatypical_Carcinoma
C510-C512,C518, C529|Vagina|809|Basal_Cell_Carcinoma|8097/3|Skin_Nodular_Basal_Cell_Carcinoma
C510-C512,C518, C529|Vagina|809|Basal_Cell_Carcinoma|8098/3|Skin_Adenoid_Basal_Cell_Carcinoma
C510-C512,C518, C529|Vagina|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C510-C512,C518, C529|Vagina|811|Pilomatrical_Carcinoma|8110/3|Pilomatrical_Carcinoma
C510-C512,C518, C529|Vagina|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C510-C512,C518, C529|Vagina|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C510-C512,C518, C529|Vagina|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C510-C512,C518, C529|Vagina|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C510-C512,C518, C529|Vagina|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C510-C512,C518, C529|Vagina|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C510-C512,C518, C529|Vagina|813|Carcinoma|8130/2|Carcinoma
C510-C512,C518, C529|Vagina|813|Carcinoma|8130/3|Carcinoma
C510-C512,C518, C529|Vagina|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8140/3|Adenocarcinoma
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C510-C512,C518, C529|Vagina|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C510-C512,C518, C529|Vagina|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C510-C512,C518, C529|Vagina|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C510-C512,C518, C529|Vagina|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C510-C512,C518, C529|Vagina|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C510-C512,C518, C529|Vagina|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C510-C512,C518, C529|Vagina|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C510-C512,C518, C529|Vagina|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C510-C512,C518, C529|Vagina|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C510-C512,C518, C529|Vagina|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C510-C512,C518, C529|Vagina|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C510-C512,C518, C529|Vagina|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C510-C512,C518, C529|Vagina|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C510-C512,C518, C529|Vagina|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C510-C512,C518, C529|Vagina|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C510-C512,C518, C529|Vagina|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C510-C512,C518, C529|Vagina|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C510-C512,C518, C529|Vagina|848|Mucinous_Adenocarcinoma|8482/3|Adenocarcinoma__Endocervical_Type
C510-C512,C518, C529|Vagina|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C510-C512,C518, C529|Vagina|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C510-C512,C518, C529|Vagina|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C510-C512,C518, C529|Vagina|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C510-C512,C518, C529|Vagina|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C510-C512,C518, C529|Vagina|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C510-C512,C518, C529|Vagina|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C510-C512,C518, C529|Vagina|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C510-C512,C518, C529|Vagina|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C510-C512,C518, C529|Vagina|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C510-C512,C518, C529|Vagina|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C510-C512,C518, C529|Vagina|872|Melanoma|8720/3|Melanoma
C510-C512,C518, C529|Vagina|872|Melanoma|8721/3|Nodular_Melanoma
C510-C512,C518, C529|Vagina|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C510-C512,C518, C529|Vagina|872|Melanoma|8723/3|Regressing_Melanoma
C510-C512,C518, C529|Vagina|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C510-C512,C518, C529|Vagina|874|Nevus|8740/3|Melanoma_In_Junctional_Nevus
C510-C512,C518, C529|Vagina|874|Nevus|8741/2|Precancerous_Melanosis
C510-C512,C518, C529|Vagina|874|Nevus|8741/3|Melanoma
C510-C512,C518, C529|Vagina|874|Nevus|8742/2|Lentigo_Maligna
C510-C512,C518, C529|Vagina|874|Nevus|8742/3|Lentigo_Maligna_Melanoma
C510-C512,C518, C529|Vagina|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C510-C512,C518, C529|Vagina|874|Nevus|8745/3|Desmoplastic_Melanoma
C510-C512,C518, C529|Vagina|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C510-C512,C518, C529|Vagina|876|Nevus|8761/3|Giant_Congenital_Nevus
C510-C512,C518, C529|Vagina|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C510-C512,C518, C529|Vagina|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C510-C512,C518, C529|Vagina|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8800/3|Sarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C510-C512,C518, C529|Vagina|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C510-C512,C518, C529|Vagina|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C510-C512,C518, C529|Vagina|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C510-C512,C518, C529|Vagina|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C510-C512,C518, C529|Vagina|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C510-C512,C518, C529|Vagina|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C510-C512,C518, C529|Vagina|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C510-C512,C518, C529|Vagina|882|Sarcoma|8825/3|Sarcoma
C510-C512,C518, C529|Vagina|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C510-C512,C518, C529|Vagina|883|Benign_Fibrous_Histiocytoma|8832/3|Dermatofibrosarcoma_Protuberans
C510-C512,C518, C529|Vagina|885|Liposarcoma|8850/3|Liposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C510-C512,C518, C529|Vagina|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8855/3|Liposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C510-C512,C518, C529|Vagina|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C510-C512,C518, C529|Vagina|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C510-C512,C518, C529|Vagina|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C510-C512,C518, C529|Vagina|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C510-C512,C518, C529|Vagina|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C510-C512,C518, C529|Vagina|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C510-C512,C518, C529|Vagina|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C510-C512,C518, C529|Vagina|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C510-C512,C518, C529|Vagina|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C510-C512,C518, C529|Vagina|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C510-C512,C518, C529|Vagina|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C510-C512,C518, C529|Vagina|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C510-C512,C518, C529|Vagina|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C510-C512,C518, C529|Vagina|898|Carcinosarcoma|8980/3|Carcinosarcoma
C510-C512,C518, C529|Vagina|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C510-C512,C518, C529|Vagina|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C510-C512,C518, C529|Vagina|911|Mesonephroma|9110/3|Mesonephroma
C510-C512,C518, C529|Vagina|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C510-C512,C518, C529|Vagina|959|Lymphoma|9590/3|Lymphoma
C510-C512,C518, C529|Vagina|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|959|Lymphoma|9597/3|Crosti_s_Disease
C510-C512,C518, C529|Vagina|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C510-C512,C518, C529|Vagina|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C510-C512,C518, C529|Vagina|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C510-C512,C518, C529|Vagina|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C510-C512,C518, C529|Vagina|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C510-C512,C518, C529|Vagina|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C510-C512,C518, C529|Vagina|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C510-C512,C518, C529|Vagina|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C510-C512,C518, C529|Vagina|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C510-C512,C518, C529|Vagina|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C510-C512,C518, C529|Vagina|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C510-C512,C518, C529|Vagina|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C510-C512,C518, C529|Vagina|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C510-C512,C518, C529|Vagina|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C510-C512,C518, C529|Vagina|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C510-C512,C518, C529|Vagina|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C510-C512,C518, C529|Vagina|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C510-C512,C518, C529|Vagina|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C510-C512,C518, C529|Vagina|970|T_Cell_Lymphoma|9700/3|Mycosis_Fungoides
C510-C512,C518, C529|Vagina|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C510-C512,C518, C529|Vagina|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C510-C512,C518, C529|Vagina|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C510-C512,C518, C529|Vagina|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C510-C512,C518, C529|Vagina|970|T_Cell_Lymphoma|9709/3|Cutaneous_T_Cell_Non_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C510-C512,C518, C529|Vagina|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C510-C512,C518, C529|Vagina|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C510-C512,C518, C529|Vagina|971|Adult_Non_Hodgkin_Lymphoma|9718/3|C_ALCL
C510-C512,C518, C529|Vagina|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C510-C512,C518, C529|Vagina|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C510-C512,C518, C529|Vagina|972|Lymphoblastic_Lymphoma|9725/3|Hydroa_Vacciniforme_Like_Lymphoma
C510-C512,C518, C529|Vagina|972|Lymphoblastic_Lymphoma|9726/3|T_Cell_Lymphoma
C510-C512,C518, C529|Vagina|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C510-C512,C518, C529|Vagina|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C510-C512,C518, C529|Vagina|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9731/3|Plasmacytoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C510-C512,C518, C529|Vagina|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C510-C512,C518, C529|Vagina|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C510-C512,C518, C529|Vagina|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C510-C512,C518, C529|Vagina|975|Neoplasm|9750/3|Malignant_Histiocytosis
C510-C512,C518, C529|Vagina|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C510-C512,C518, C529|Vagina|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C510-C512,C518, C529|Vagina|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C510-C512,C518, C529|Vagina|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C510-C512,C518, C529|Vagina|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C510-C512,C518, C529|Vagina|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C510-C512,C518, C529|Vagina|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C510-C512,C518, C529|Vagina|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C510-C512,C518, C529|Vagina|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C510-C512,C518, C529|Vagina|981|Neoplasm|9812/3|Lymphoma
C510-C512,C518, C529|Vagina|981|Neoplasm|9813/3|Lymphoma
C510-C512,C518, C529|Vagina|981|Neoplasm|9814/3|Lymphoma
C510-C512,C518, C529|Vagina|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C510-C512,C518, C529|Vagina|981|Neoplasm|9816/3|Hypodiploid_ALL
C510-C512,C518, C529|Vagina|981|Neoplasm|9817/3|Lymphoma
C510-C512,C518, C529|Vagina|981|Neoplasm|9818/3|Lymphoma
C510-C512,C518, C529|Vagina|981|Neoplasm|9819/3|Leukemia__B_Cell
C510-C512,C518, C529|Vagina|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C510-C512,C518, C529|Vagina|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C510-C512,C518, C529|Vagina|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C510-C512,C518, C529|Vagina|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C510-C512,C518, C529|Vagina|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C510-C512,C518, C529|Vagina|997|Neoplasm|9971/3|Polymorphic_PTLD
C510-C512,C518, C529|Vagina|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C519|Vulva|800|Neoplasm|8000/3|Malignant_Neoplasm
C519|Vulva|800|Neoplasm|8001/3|Malignant_Cell
C519|Vulva|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C519|Vulva|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C519|Vulva|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C519|Vulva|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C519|Vulva|801|Carcinoma|8010/2|In_Situ_Cancer
C519|Vulva|801|Carcinoma|8010/3|Carcinoma
C519|Vulva|801|Carcinoma|8011/3|Malignant_Epithelioma
C519|Vulva|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C519|Vulva|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C519|Vulva|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C519|Vulva|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C519|Vulva|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C519|Vulva|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C519|Vulva|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C519|Vulva|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C519|Vulva|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C519|Vulva|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C519|Vulva|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C519|Vulva|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C519|Vulva|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8071/2|Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C519|Vulva|807|Squamous_Cell_Carcinoma|8077/2|Intraepithelial_Neoplasia
C519|Vulva|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C519|Vulva|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C519|Vulva|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C519|Vulva|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C519|Vulva|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C519|Vulva|809|Basal_Cell_Carcinoma|8090/3|Basal_Cell_Carcinoma
C519|Vulva|809|Basal_Cell_Carcinoma|8091/3|Superficial_Basal_Cell_Carcinoma
C519|Vulva|809|Basal_Cell_Carcinoma|8092/3|Skin_Infiltrating_Basal_Cell_Carcinoma
C519|Vulva|809|Basal_Cell_Carcinoma|8093/3|Fibroepithelioma_Of_Pinkus
C519|Vulva|809|Basal_Cell_Carcinoma|8094/3|Skin_Basosquamous_Cell_Carcinoma
C519|Vulva|809|Basal_Cell_Carcinoma|8095/3|Skin_Metatypical_Carcinoma
C519|Vulva|809|Basal_Cell_Carcinoma|8097/3|Skin_Nodular_Basal_Cell_Carcinoma
C519|Vulva|809|Basal_Cell_Carcinoma|8098/3|Skin_Adenoid_Basal_Cell_Carcinoma
C519|Vulva|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C519|Vulva|811|Pilomatrical_Carcinoma|8110/3|Pilomatrical_Carcinoma
C519|Vulva|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C519|Vulva|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C519|Vulva|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C519|Vulva|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C519|Vulva|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C519|Vulva|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C519|Vulva|813|Carcinoma|8130/2|Carcinoma
C519|Vulva|813|Carcinoma|8130/3|Carcinoma
C519|Vulva|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C519|Vulva|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C519|Vulva|814|Adenocarcinoma|8140/3|Adenocarcinoma
C519|Vulva|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C519|Vulva|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C519|Vulva|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C519|Vulva|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C519|Vulva|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C519|Vulva|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C519|Vulva|824|Atypical_Carcinoid_Tumor|8247/3|Merkel_Cell_Carcinoma
C519|Vulva|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C519|Vulva|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C519|Vulva|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C519|Vulva|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C519|Vulva|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C519|Vulva|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C519|Vulva|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C519|Vulva|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C519|Vulva|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C519|Vulva|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C519|Vulva|839|Adnexal_Carcinoma|8390/3|Adnexal_Carcinoma
C519|Vulva|840|Sweat_Gland_Adenocarcinoma|8400/3|Sweat_Gland_Adenocarcinoma
C519|Vulva|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C519|Vulva|841|Eccrine_Adenocarcinoma|8410/3|Sebaceous_Adenocarcinoma
C519|Vulva|841|Eccrine_Adenocarcinoma|8413/3|Eccrine_Adenocarcinoma
C519|Vulva|842|Ceruminous_Adenocarcinoma|8420/3|Ceruminous_Adenocarcinoma
C519|Vulva|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C519|Vulva|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C519|Vulva|848|Mucinous_Adenocarcinoma|8482/3|Adenocarcinoma__Endocervical_Type
C519|Vulva|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C519|Vulva|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C519|Vulva|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C519|Vulva|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C519|Vulva|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C519|Vulva|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C519|Vulva|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C519|Vulva|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C519|Vulva|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C519|Vulva|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C519|Vulva|872|Melanoma|8720/3|Melanoma
C519|Vulva|872|Melanoma|8721/3|Nodular_Melanoma
C519|Vulva|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C519|Vulva|872|Melanoma|8723/3|Regressing_Melanoma
C519|Vulva|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C519|Vulva|874|Nevus|8740/3|Melanoma_In_Junctional_Nevus
C519|Vulva|874|Nevus|8741/2|Precancerous_Melanosis
C519|Vulva|874|Nevus|8741/3|Melanoma
C519|Vulva|874|Nevus|8742/2|Lentigo_Maligna
C519|Vulva|874|Nevus|8742/3|Lentigo_Maligna_Melanoma
C519|Vulva|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C519|Vulva|874|Nevus|8745/3|Desmoplastic_Melanoma
C519|Vulva|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C519|Vulva|876|Nevus|8761/3|Giant_Congenital_Nevus
C519|Vulva|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C519|Vulva|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C519|Vulva|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C519|Vulva|878|Melanoma_Arising_From_Blue_Nevus|8780/3|Melanoma_Arising_From_Blue_Nevus
C519|Vulva|880|Sarcoma|8800/3|Sarcoma
C519|Vulva|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C519|Vulva|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C519|Vulva|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C519|Vulva|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C519|Vulva|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C519|Vulva|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C519|Vulva|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C519|Vulva|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C519|Vulva|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C519|Vulva|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C519|Vulva|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C519|Vulva|882|Sarcoma|8825/3|Sarcoma
C519|Vulva|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C519|Vulva|883|Benign_Fibrous_Histiocytoma|8832/3|Dermatofibrosarcoma_Protuberans
C519|Vulva|885|Liposarcoma|8850/3|Liposarcoma
C519|Vulva|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C519|Vulva|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C519|Vulva|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C519|Vulva|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C519|Vulva|885|Liposarcoma|8855/3|Liposarcoma
C519|Vulva|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C519|Vulva|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C519|Vulva|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C519|Vulva|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C519|Vulva|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C519|Vulva|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C519|Vulva|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C519|Vulva|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C519|Vulva|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C519|Vulva|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C519|Vulva|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C519|Vulva|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C519|Vulva|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C519|Vulva|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C519|Vulva|898|Carcinosarcoma|8980/3|Carcinosarcoma
C519|Vulva|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C519|Vulva|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C519|Vulva|911|Mesonephroma|9110/3|Mesonephroma
C519|Vulva|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C519|Vulva|959|Lymphoma|9590/3|Lymphoma
C519|Vulva|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C519|Vulva|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C519|Vulva|959|Lymphoma|9597/3|Crosti_s_Disease
C519|Vulva|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C519|Vulva|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C519|Vulva|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C519|Vulva|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C519|Vulva|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C519|Vulva|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C519|Vulva|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C519|Vulva|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C519|Vulva|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C519|Vulva|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C519|Vulva|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C519|Vulva|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C519|Vulva|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C519|Vulva|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C519|Vulva|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C519|Vulva|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C519|Vulva|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C519|Vulva|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C519|Vulva|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C519|Vulva|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C519|Vulva|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C519|Vulva|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C519|Vulva|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C519|Vulva|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C519|Vulva|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C519|Vulva|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C519|Vulva|970|T_Cell_Lymphoma|9700/3|Mycosis_Fungoides
C519|Vulva|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C519|Vulva|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C519|Vulva|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C519|Vulva|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C519|Vulva|970|T_Cell_Lymphoma|9709/3|Cutaneous_T_Cell_Non_Hodgkin_Lymphoma
C519|Vulva|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C519|Vulva|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C519|Vulva|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C519|Vulva|971|Adult_Non_Hodgkin_Lymphoma|9718/3|C_ALCL
C519|Vulva|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C519|Vulva|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C519|Vulva|972|Lymphoblastic_Lymphoma|9725/3|Hydroa_Vacciniforme_Like_Lymphoma
C519|Vulva|972|Lymphoblastic_Lymphoma|9726/3|T_Cell_Lymphoma
C519|Vulva|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C519|Vulva|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C519|Vulva|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C519|Vulva|973|Plasmacytoma|9731/3|Plasmacytoma
C519|Vulva|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C519|Vulva|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C519|Vulva|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C519|Vulva|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C519|Vulva|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C519|Vulva|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C519|Vulva|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C519|Vulva|975|Neoplasm|9750/3|Malignant_Histiocytosis
C519|Vulva|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C519|Vulva|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C519|Vulva|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C519|Vulva|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C519|Vulva|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C519|Vulva|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C519|Vulva|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C519|Vulva|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C519|Vulva|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C519|Vulva|981|Neoplasm|9812/3|Lymphoma
C519|Vulva|981|Neoplasm|9813/3|Lymphoma
C519|Vulva|981|Neoplasm|9814/3|Lymphoma
C519|Vulva|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C519|Vulva|981|Neoplasm|9816/3|Hypodiploid_ALL
C519|Vulva|981|Neoplasm|9817/3|Lymphoma
C519|Vulva|981|Neoplasm|9818/3|Lymphoma
C519|Vulva|981|Neoplasm|9819/3|Leukemia__B_Cell
C519|Vulva|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C519|Vulva|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C519|Vulva|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C519|Vulva|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C519|Vulva|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C519|Vulva|997|Neoplasm|9971/3|Polymorphic_PTLD
C519|Vulva|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C530-C531,C538-C539|Cervix_Uteri|800|Neoplasm|8000/3|Malignant_Neoplasm
C530-C531,C538-C539|Cervix_Uteri|800|Neoplasm|8001/3|Malignant_Cell
C530-C531,C538-C539|Cervix_Uteri|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C530-C531,C538-C539|Cervix_Uteri|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C530-C531,C538-C539|Cervix_Uteri|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C530-C531,C538-C539|Cervix_Uteri|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C530-C531,C538-C539|Cervix_Uteri|801|Carcinoma|8010/2|In_Situ_Cancer
C530-C531,C538-C539|Cervix_Uteri|801|Carcinoma|8010/3|Carcinoma
C530-C531,C538-C539|Cervix_Uteri|801|Carcinoma|8011/3|Malignant_Epithelioma
C530-C531,C538-C539|Cervix_Uteri|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C530-C531,C538-C539|Cervix_Uteri|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C530-C531,C538-C539|Cervix_Uteri|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C530-C531,C538-C539|Cervix_Uteri|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8071/2|Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8072/2|Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8077/2|Intraepithelial_Neoplasia
C530-C531,C538-C539|Cervix_Uteri|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C530-C531,C538-C539|Cervix_Uteri|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|809|Basal_Cell_Carcinoma|8098/3|Skin_Adenoid_Basal_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C530-C531,C538-C539|Cervix_Uteri|814|Adenocarcinoma|8140/3|Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C530-C531,C538-C539|Cervix_Uteri|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C530-C531,C538-C539|Cervix_Uteri|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C530-C531,C538-C539|Cervix_Uteri|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C530-C531,C538-C539|Cervix_Uteri|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C530-C531,C538-C539|Cervix_Uteri|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C530-C531,C538-C539|Cervix_Uteri|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C530-C531,C538-C539|Cervix_Uteri|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|838|Carcinoma__Endometrioid|8384/3|Adenocarcinoma__Endocervical_Type
C530-C531,C538-C539|Cervix_Uteri|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|848|Mucinous_Adenocarcinoma|8482/3|Adenocarcinoma__Endocervical_Type
C530-C531,C538-C539|Cervix_Uteri|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C530-C531,C538-C539|Cervix_Uteri|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C530-C531,C538-C539|Cervix_Uteri|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C530-C531,C538-C539|Cervix_Uteri|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C530-C531,C538-C539|Cervix_Uteri|880|Sarcoma|8800/3|Sarcoma
C530-C531,C538-C539|Cervix_Uteri|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C530-C531,C538-C539|Cervix_Uteri|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C530-C531,C538-C539|Cervix_Uteri|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C530-C531,C538-C539|Cervix_Uteri|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C530-C531,C538-C539|Cervix_Uteri|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C530-C531,C538-C539|Cervix_Uteri|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C530-C531,C538-C539|Cervix_Uteri|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C530-C531,C538-C539|Cervix_Uteri|882|Sarcoma|8825/3|Sarcoma
C530-C531,C538-C539|Cervix_Uteri|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C530-C531,C538-C539|Cervix_Uteri|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C530-C531,C538-C539|Cervix_Uteri|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C530-C531,C538-C539|Cervix_Uteri|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C530-C531,C538-C539|Cervix_Uteri|898|Carcinosarcoma|8980/3|Carcinosarcoma
C530-C531,C538-C539|Cervix_Uteri|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C530-C531,C538-C539|Cervix_Uteri|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C530-C531,C538-C539|Cervix_Uteri|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C530-C531,C538-C539|Cervix_Uteri|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C530-C531,C538-C539|Cervix_Uteri|911|Mesonephroma|9110/3|Mesonephroma
C530-C531,C538-C539|Cervix_Uteri|959|Lymphoma|9590/3|Lymphoma
C530-C531,C538-C539|Cervix_Uteri|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C530-C531,C538-C539|Cervix_Uteri|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C530-C531,C538-C539|Cervix_Uteri|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C530-C531,C538-C539|Cervix_Uteri|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C530-C531,C538-C539|Cervix_Uteri|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C530-C531,C538-C539|Cervix_Uteri|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C530-C531,C538-C539|Cervix_Uteri|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C530-C531,C538-C539|Cervix_Uteri|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C530-C531,C538-C539|Cervix_Uteri|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C530-C531,C538-C539|Cervix_Uteri|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C530-C531,C538-C539|Cervix_Uteri|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C530-C531,C538-C539|Cervix_Uteri|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C530-C531,C538-C539|Cervix_Uteri|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C530-C531,C538-C539|Cervix_Uteri|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|973|Plasmacytoma|9731/3|Plasmacytoma
C530-C531,C538-C539|Cervix_Uteri|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C530-C531,C538-C539|Cervix_Uteri|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C530-C531,C538-C539|Cervix_Uteri|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C530-C531,C538-C539|Cervix_Uteri|975|Neoplasm|9750/3|Malignant_Histiocytosis
C530-C531,C538-C539|Cervix_Uteri|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C530-C531,C538-C539|Cervix_Uteri|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C530-C531,C538-C539|Cervix_Uteri|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C530-C531,C538-C539|Cervix_Uteri|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C530-C531,C538-C539|Cervix_Uteri|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9812/3|Lymphoma
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9813/3|Lymphoma
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9814/3|Lymphoma
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9816/3|Hypodiploid_ALL
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9817/3|Lymphoma
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9818/3|Lymphoma
C530-C531,C538-C539|Cervix_Uteri|981|Neoplasm|9819/3|Leukemia__B_Cell
C530-C531,C538-C539|Cervix_Uteri|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C530-C531,C538-C539|Cervix_Uteri|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C530-C531,C538-C539|Cervix_Uteri|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C530-C531,C538-C539|Cervix_Uteri|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C530-C531,C538-C539|Cervix_Uteri|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C530-C531,C538-C539|Cervix_Uteri|997|Neoplasm|9971/3|Polymorphic_PTLD
C530-C531,C538-C539|Cervix_Uteri|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C540-C543,C548-C549|Corpus_Uteri|800|Neoplasm|8000/3|Malignant_Neoplasm
C540-C543,C548-C549|Corpus_Uteri|800|Neoplasm|8001/3|Malignant_Cell
C540-C543,C548-C549|Corpus_Uteri|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C540-C543,C548-C549|Corpus_Uteri|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C540-C543,C548-C549|Corpus_Uteri|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C540-C543,C548-C549|Corpus_Uteri|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C540-C543,C548-C549|Corpus_Uteri|801|Carcinoma|8010/2|In_Situ_Cancer
C540-C543,C548-C549|Corpus_Uteri|801|Carcinoma|8010/3|Carcinoma
C540-C543,C548-C549|Corpus_Uteri|801|Carcinoma|8011/3|Malignant_Epithelioma
C540-C543,C548-C549|Corpus_Uteri|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C540-C543,C548-C549|Corpus_Uteri|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C540-C543,C548-C549|Corpus_Uteri|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C540-C543,C548-C549|Corpus_Uteri|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C540-C543,C548-C549|Corpus_Uteri|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|813|Carcinoma|8130/2|Carcinoma
C540-C543,C548-C549|Corpus_Uteri|813|Carcinoma|8130/3|Carcinoma
C540-C543,C548-C549|Corpus_Uteri|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C540-C543,C548-C549|Corpus_Uteri|814|Adenocarcinoma|8140/3|Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C540-C543,C548-C549|Corpus_Uteri|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C540-C543,C548-C549|Corpus_Uteri|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C540-C543,C548-C549|Corpus_Uteri|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C540-C543,C548-C549|Corpus_Uteri|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C540-C543,C548-C549|Corpus_Uteri|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C540-C543,C548-C549|Corpus_Uteri|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C540-C543,C548-C549|Corpus_Uteri|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C540-C543,C548-C549|Corpus_Uteri|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C540-C543,C548-C549|Corpus_Uteri|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C540-C543,C548-C549|Corpus_Uteri|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|838|Carcinoma__Endometrioid|8380/2|Atypical_Endometrial_Hyperplasia
C540-C543,C548-C549|Corpus_Uteri|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C540-C543,C548-C549|Corpus_Uteri|838|Carcinoma__Endometrioid|8381/3|Endometrioid_Adenofibroma__Malignant
C540-C543,C548-C549|Corpus_Uteri|838|Carcinoma__Endometrioid|8382/3|Carcinoma__Endometrioid
C540-C543,C548-C549|Corpus_Uteri|838|Carcinoma__Endometrioid|8383/3|Carcinoma__Endometrioid
C540-C543,C548-C549|Corpus_Uteri|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|844|Cystadenocarcinoma|8441/2|Serous_Tubal_Intraepithelial_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|844|Cystadenocarcinoma|8441/3|Serous_Cystadenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|846|Papillary_Serous_Cystadenocarcinoma|8460/3|Papillary_Serous_Cystadenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|846|Papillary_Serous_Cystadenocarcinoma|8461/3|Serous_Surface_Papillary_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|848|Mucinous_Adenocarcinoma|8482/3|Adenocarcinoma__Endocervical_Type
C540-C543,C548-C549|Corpus_Uteri|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C540-C543,C548-C549|Corpus_Uteri|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C540-C543,C548-C549|Corpus_Uteri|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C540-C543,C548-C549|Corpus_Uteri|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C540-C543,C548-C549|Corpus_Uteri|880|Sarcoma|8800/3|Sarcoma
C540-C543,C548-C549|Corpus_Uteri|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C540-C543,C548-C549|Corpus_Uteri|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C540-C543,C548-C549|Corpus_Uteri|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C540-C543,C548-C549|Corpus_Uteri|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C540-C543,C548-C549|Corpus_Uteri|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C540-C543,C548-C549|Corpus_Uteri|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C540-C543,C548-C549|Corpus_Uteri|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C540-C543,C548-C549|Corpus_Uteri|882|Sarcoma|8825/3|Sarcoma
C540-C543,C548-C549|Corpus_Uteri|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C540-C543,C548-C549|Corpus_Uteri|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C540-C543,C548-C549|Corpus_Uteri|893|Stromal_Sarcoma|8930/3|Endometrial_Stromal_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|893|Stromal_Sarcoma|8931/3|Low_Grade_Endometrioid_Stromal_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|893|Stromal_Sarcoma|8933/3|Adenosarcoma
C540-C543,C548-C549|Corpus_Uteri|893|Stromal_Sarcoma|8934/3|Carcinofibroma
C540-C543,C548-C549|Corpus_Uteri|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C540-C543,C548-C549|Corpus_Uteri|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C540-C543,C548-C549|Corpus_Uteri|898|Carcinosarcoma|8980/3|Carcinosarcoma
C540-C543,C548-C549|Corpus_Uteri|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C540-C543,C548-C549|Corpus_Uteri|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C540-C543,C548-C549|Corpus_Uteri|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C540-C543,C548-C549|Corpus_Uteri|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C540-C543,C548-C549|Corpus_Uteri|911|Mesonephroma|9110/3|Mesonephroma
C540-C543,C548-C549|Corpus_Uteri|959|Lymphoma|9590/3|Lymphoma
C540-C543,C548-C549|Corpus_Uteri|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C540-C543,C548-C549|Corpus_Uteri|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C540-C543,C548-C549|Corpus_Uteri|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C540-C543,C548-C549|Corpus_Uteri|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C540-C543,C548-C549|Corpus_Uteri|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C540-C543,C548-C549|Corpus_Uteri|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C540-C543,C548-C549|Corpus_Uteri|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C540-C543,C548-C549|Corpus_Uteri|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C540-C543,C548-C549|Corpus_Uteri|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C540-C543,C548-C549|Corpus_Uteri|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C540-C543,C548-C549|Corpus_Uteri|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C540-C543,C548-C549|Corpus_Uteri|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C540-C543,C548-C549|Corpus_Uteri|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C540-C543,C548-C549|Corpus_Uteri|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|973|Plasmacytoma|9731/3|Plasmacytoma
C540-C543,C548-C549|Corpus_Uteri|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C540-C543,C548-C549|Corpus_Uteri|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C540-C543,C548-C549|Corpus_Uteri|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C540-C543,C548-C549|Corpus_Uteri|975|Neoplasm|9750/3|Malignant_Histiocytosis
C540-C543,C548-C549|Corpus_Uteri|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C540-C543,C548-C549|Corpus_Uteri|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C540-C543,C548-C549|Corpus_Uteri|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C540-C543,C548-C549|Corpus_Uteri|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C540-C543,C548-C549|Corpus_Uteri|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9812/3|Lymphoma
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9813/3|Lymphoma
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9814/3|Lymphoma
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9816/3|Hypodiploid_ALL
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9817/3|Lymphoma
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9818/3|Lymphoma
C540-C543,C548-C549|Corpus_Uteri|981|Neoplasm|9819/3|Leukemia__B_Cell
C540-C543,C548-C549|Corpus_Uteri|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C540-C543,C548-C549|Corpus_Uteri|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C540-C543,C548-C549|Corpus_Uteri|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C540-C543,C548-C549|Corpus_Uteri|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C540-C543,C548-C549|Corpus_Uteri|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C540-C543,C548-C549|Corpus_Uteri|997|Neoplasm|9971/3|Polymorphic_PTLD
C540-C543,C548-C549|Corpus_Uteri|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C559|Uterus|800|Neoplasm|8000/3|Malignant_Neoplasm
C559|Uterus|800|Neoplasm|8001/3|Malignant_Cell
C559|Uterus|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C559|Uterus|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C559|Uterus|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C559|Uterus|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C559|Uterus|801|Carcinoma|8010/2|In_Situ_Cancer
C559|Uterus|801|Carcinoma|8010/3|Carcinoma
C559|Uterus|801|Carcinoma|8011/3|Malignant_Epithelioma
C559|Uterus|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C559|Uterus|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C559|Uterus|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C559|Uterus|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C559|Uterus|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C559|Uterus|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C559|Uterus|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C559|Uterus|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C559|Uterus|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C559|Uterus|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C559|Uterus|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C559|Uterus|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C559|Uterus|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C559|Uterus|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C559|Uterus|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C559|Uterus|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C559|Uterus|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C559|Uterus|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C559|Uterus|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C559|Uterus|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C559|Uterus|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C559|Uterus|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C559|Uterus|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C559|Uterus|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C559|Uterus|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C559|Uterus|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C559|Uterus|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C559|Uterus|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C559|Uterus|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C559|Uterus|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C559|Uterus|813|Carcinoma|8130/2|Carcinoma
C559|Uterus|813|Carcinoma|8130/3|Carcinoma
C559|Uterus|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C559|Uterus|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C559|Uterus|814|Adenocarcinoma|8140/3|Adenocarcinoma
C559|Uterus|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C559|Uterus|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C559|Uterus|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C559|Uterus|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C559|Uterus|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C559|Uterus|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C559|Uterus|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C559|Uterus|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C559|Uterus|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C559|Uterus|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C559|Uterus|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C559|Uterus|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C559|Uterus|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C559|Uterus|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C559|Uterus|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C559|Uterus|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C559|Uterus|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C559|Uterus|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C559|Uterus|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C559|Uterus|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C559|Uterus|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C559|Uterus|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C559|Uterus|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C559|Uterus|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C559|Uterus|844|Cystadenocarcinoma|8441/2|Serous_Tubal_Intraepithelial_Carcinoma
C559|Uterus|844|Cystadenocarcinoma|8441/3|Serous_Cystadenocarcinoma
C559|Uterus|846|Papillary_Serous_Cystadenocarcinoma|8460/3|Papillary_Serous_Cystadenocarcinoma
C559|Uterus|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C559|Uterus|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C559|Uterus|848|Mucinous_Adenocarcinoma|8482/3|Adenocarcinoma__Endocervical_Type
C559|Uterus|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C559|Uterus|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C559|Uterus|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C559|Uterus|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C559|Uterus|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C559|Uterus|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C559|Uterus|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C559|Uterus|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C559|Uterus|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C559|Uterus|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C559|Uterus|880|Sarcoma|8800/3|Sarcoma
C559|Uterus|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C559|Uterus|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C559|Uterus|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C559|Uterus|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C559|Uterus|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C559|Uterus|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C559|Uterus|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C559|Uterus|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C559|Uterus|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C559|Uterus|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C559|Uterus|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C559|Uterus|882|Sarcoma|8825/3|Sarcoma
C559|Uterus|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C559|Uterus|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C559|Uterus|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C559|Uterus|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C559|Uterus|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C559|Uterus|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C559|Uterus|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C559|Uterus|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C559|Uterus|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C559|Uterus|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C559|Uterus|893|Stromal_Sarcoma|8930/3|Endometrial_Stromal_Sarcoma
C559|Uterus|893|Stromal_Sarcoma|8931/3|Low_Grade_Endometrioid_Stromal_Sarcoma
C559|Uterus|893|Stromal_Sarcoma|8934/3|Carcinofibroma
C559|Uterus|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C559|Uterus|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C559|Uterus|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C559|Uterus|898|Carcinosarcoma|8980/3|Carcinosarcoma
C559|Uterus|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C559|Uterus|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C559|Uterus|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C559|Uterus|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C559|Uterus|911|Mesonephroma|9110/3|Mesonephroma
C559|Uterus|959|Lymphoma|9590/3|Lymphoma
C559|Uterus|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C559|Uterus|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C559|Uterus|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C559|Uterus|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C559|Uterus|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C559|Uterus|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C559|Uterus|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C559|Uterus|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C559|Uterus|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C559|Uterus|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C559|Uterus|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C559|Uterus|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C559|Uterus|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C559|Uterus|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C559|Uterus|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C559|Uterus|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C559|Uterus|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C559|Uterus|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C559|Uterus|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C559|Uterus|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C559|Uterus|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C559|Uterus|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C559|Uterus|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C559|Uterus|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C559|Uterus|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C559|Uterus|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C559|Uterus|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C559|Uterus|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C559|Uterus|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C559|Uterus|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C559|Uterus|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C559|Uterus|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C559|Uterus|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C559|Uterus|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C559|Uterus|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C559|Uterus|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C559|Uterus|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C559|Uterus|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C559|Uterus|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C559|Uterus|973|Plasmacytoma|9731/3|Plasmacytoma
C559|Uterus|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C559|Uterus|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C559|Uterus|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C559|Uterus|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C559|Uterus|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C559|Uterus|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C559|Uterus|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C559|Uterus|975|Neoplasm|9750/3|Malignant_Histiocytosis
C559|Uterus|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C559|Uterus|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C559|Uterus|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C559|Uterus|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C559|Uterus|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C559|Uterus|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C559|Uterus|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C559|Uterus|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C559|Uterus|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C559|Uterus|981|Neoplasm|9812/3|Lymphoma
C559|Uterus|981|Neoplasm|9813/3|Lymphoma
C559|Uterus|981|Neoplasm|9814/3|Lymphoma
C559|Uterus|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C559|Uterus|981|Neoplasm|9816/3|Hypodiploid_ALL
C559|Uterus|981|Neoplasm|9817/3|Lymphoma
C559|Uterus|981|Neoplasm|9818/3|Lymphoma
C559|Uterus|981|Neoplasm|9819/3|Leukemia__B_Cell
C559|Uterus|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C559|Uterus|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C559|Uterus|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C559|Uterus|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C559|Uterus|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C559|Uterus|997|Neoplasm|9971/3|Polymorphic_PTLD
C559|Uterus|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C569|Ovary|800|Neoplasm|8000/3|Malignant_Neoplasm
C569|Ovary|800|Neoplasm|8001/3|Malignant_Cell
C569|Ovary|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C569|Ovary|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C569|Ovary|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C569|Ovary|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C569|Ovary|801|Carcinoma|8010/2|In_Situ_Cancer
C569|Ovary|801|Carcinoma|8010/3|Carcinoma
C569|Ovary|801|Carcinoma|8011/3|Malignant_Epithelioma
C569|Ovary|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C569|Ovary|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C569|Ovary|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C569|Ovary|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C569|Ovary|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C569|Ovary|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C569|Ovary|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C569|Ovary|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C569|Ovary|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C569|Ovary|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C569|Ovary|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C569|Ovary|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C569|Ovary|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C569|Ovary|804|Small_Cell_Carcinoma|8041/3|Ovarian_Small_Cell_Carcinoma
C569|Ovary|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C569|Ovary|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C569|Ovary|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C569|Ovary|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C569|Ovary|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C569|Ovary|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C569|Ovary|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C569|Ovary|814|Adenocarcinoma|8140/3|Adenocarcinoma
C569|Ovary|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C569|Ovary|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C569|Ovary|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C569|Ovary|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C569|Ovary|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C569|Ovary|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C569|Ovary|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C569|Ovary|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C569|Ovary|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C569|Ovary|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C569|Ovary|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C569|Ovary|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C569|Ovary|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C569|Ovary|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C569|Ovary|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C569|Ovary|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C569|Ovary|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C569|Ovary|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C569|Ovary|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C569|Ovary|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C569|Ovary|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C569|Ovary|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C569|Ovary|831|Clear_Cell_Adenocarcinoma|8313/3|Clear_Cell_Adenocarcinofibroma
C569|Ovary|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C569|Ovary|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C569|Ovary|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C569|Ovary|838|Carcinoma__Endometrioid|8381/3|Endometrioid_Adenofibroma__Malignant
C569|Ovary|838|Carcinoma__Endometrioid|8382/3|Carcinoma__Endometrioid
C569|Ovary|838|Carcinoma__Endometrioid|8383/3|Carcinoma__Endometrioid
C569|Ovary|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C569|Ovary|844|Cystadenocarcinoma|8441/2|Serous_Tubal_Intraepithelial_Carcinoma
C569|Ovary|844|Cystadenocarcinoma|8441/3|Serous_Cystadenocarcinoma
C569|Ovary|844|Cystadenocarcinoma|8442/1|Serous_Cystadenoma
C569|Ovary|845|Papillary_Cystadenocarcinoma|8450/3|Papillary_Cystadenocarcinoma
C569|Ovary|845|Papillary_Cystadenocarcinoma|8451/1|Papillary_Cystadenoma
C569|Ovary|846|Papillary_Serous_Cystadenocarcinoma|8460/2|Serous_Cystadenocarcinoma
C569|Ovary|846|Papillary_Serous_Cystadenocarcinoma|8460/3|Papillary_Serous_Cystadenocarcinoma
C569|Ovary|846|Papillary_Serous_Cystadenocarcinoma|8461/3|Serous_Surface_Papillary_Carcinoma
C569|Ovary|846|Papillary_Serous_Cystadenocarcinoma|8462/1|Papillary_Cystic_Neoplasm
C569|Ovary|847|Mucinous_Cystadenocarcinoma|8470/2|Mucinous_Cystadenocarcinoma
C569|Ovary|847|Mucinous_Cystadenocarcinoma|8470/3|Mucinous_Cystadenocarcinoma
C569|Ovary|847|Mucinous_Cystadenocarcinoma|8471/3|Papillary_Mucinous_Cystadenocarcinoma
C569|Ovary|847|Mucinous_Cystadenocarcinoma|8472/1|Cystic_Neoplasm
C569|Ovary|847|Mucinous_Cystadenocarcinoma|8473/1|Papillary_Mucinous_Cystadenoma
C569|Ovary|847|Mucinous_Cystadenocarcinoma|8474/3|Carcinoma
C569|Ovary|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C569|Ovary|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C569|Ovary|848|Mucinous_Adenocarcinoma|8482/3|Adenocarcinoma__Endocervical_Type
C569|Ovary|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C569|Ovary|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C569|Ovary|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C569|Ovary|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C569|Ovary|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C569|Ovary|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C569|Ovary|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C569|Ovary|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C569|Ovary|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C569|Ovary|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C569|Ovary|859|Ovarian_Sex_Cord_Stromal_Tumor|8590/3|Ovarian_Sex_Cord_Stromal_Tumor
C569|Ovary|860|Malignant_Ovarian_Thecoma|8600/3|Malignant_Ovarian_Thecoma
C569|Ovary|862|Granulosa_Cell_Tumor|8620/3|Malignant_Granulosa_Cell_Tumor
C569|Ovary|862|Granulosa_Cell_Tumor|8621/3|Granulosa_Cell_Theca_Cell_Tumor
C569|Ovary|863|Neoplasm|8630/3|Malignant_Sertoli_Cell_Tumor
C569|Ovary|863|Neoplasm|8631/3|Sertoli_Leydig_Cell_Tumor
C569|Ovary|863|Neoplasm|8632/3|Ovarian_Gynandroblastoma
C569|Ovary|863|Neoplasm|8634/3|Sertoli_Leydig_Cell_Tumor
C569|Ovary|867|Neoplasm|8670/3|Steroid_Cell_Tumor__Malignant
C569|Ovary|880|Sarcoma|8800/3|Sarcoma
C569|Ovary|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C569|Ovary|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C569|Ovary|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C569|Ovary|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C569|Ovary|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C569|Ovary|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C569|Ovary|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C569|Ovary|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C569|Ovary|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C569|Ovary|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C569|Ovary|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C569|Ovary|882|Sarcoma|8825/3|Sarcoma
C569|Ovary|884|Myxosarcoma|8840/3|Myxosarcoma
C569|Ovary|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C569|Ovary|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C569|Ovary|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C569|Ovary|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C569|Ovary|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C569|Ovary|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C569|Ovary|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C569|Ovary|898|Carcinosarcoma|8980/3|Carcinosarcoma
C569|Ovary|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C569|Ovary|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C569|Ovary|900|Malignant_Ovarian_Brenner_Tumor|9000/3|Malignant_Ovarian_Brenner_Tumor
C569|Ovary|901|Adenocarcinofibroma|9014/3|Serous_Adenocarcinofibroma
C569|Ovary|901|Adenocarcinofibroma|9015/3|Mucinous_Adenocarcinofibroma
C569|Ovary|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C569|Ovary|906|Germ_Cell_Tumor|9064/3|Germinoma
C569|Ovary|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C569|Ovary|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C569|Ovary|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C569|Ovary|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C569|Ovary|908|Teratoma|9080/3|Immature_Teratoma
C569|Ovary|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C569|Ovary|908|Teratoma|9082/3|Immature_Teratoma
C569|Ovary|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C569|Ovary|908|Teratoma|9084/3|Teratoma
C569|Ovary|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C569|Ovary|909|Malignant_Struma_Ovarii|9090/3|Malignant_Struma_Ovarii
C569|Ovary|910|Choriocarcinoma|9100/3|Choriocarcinoma
C569|Ovary|910|Choriocarcinoma|9101/3|Choriocarcinoma
C569|Ovary|910|Choriocarcinoma|9105/3|Epithelioid_Trophoblastic_Tumor
C569|Ovary|911|Mesonephroma|9110/3|Mesonephroma
C569|Ovary|959|Lymphoma|9590/3|Lymphoma
C569|Ovary|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C569|Ovary|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C569|Ovary|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C569|Ovary|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C569|Ovary|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C569|Ovary|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C569|Ovary|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C569|Ovary|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C569|Ovary|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C569|Ovary|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C569|Ovary|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C569|Ovary|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C569|Ovary|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C569|Ovary|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C569|Ovary|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C569|Ovary|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C569|Ovary|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C569|Ovary|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C569|Ovary|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C569|Ovary|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C569|Ovary|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C569|Ovary|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C569|Ovary|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C569|Ovary|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C569|Ovary|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C569|Ovary|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C569|Ovary|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C569|Ovary|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C569|Ovary|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C569|Ovary|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C569|Ovary|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C569|Ovary|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C569|Ovary|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C569|Ovary|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C569|Ovary|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C569|Ovary|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C569|Ovary|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C569|Ovary|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C569|Ovary|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C569|Ovary|973|Plasmacytoma|9731/3|Plasmacytoma
C569|Ovary|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C569|Ovary|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C569|Ovary|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C569|Ovary|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C569|Ovary|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C569|Ovary|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C569|Ovary|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C569|Ovary|975|Neoplasm|9750/3|Malignant_Histiocytosis
C569|Ovary|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C569|Ovary|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C569|Ovary|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C569|Ovary|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C569|Ovary|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C569|Ovary|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C569|Ovary|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C569|Ovary|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C569|Ovary|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C569|Ovary|981|Neoplasm|9812/3|Lymphoma
C569|Ovary|981|Neoplasm|9813/3|Lymphoma
C569|Ovary|981|Neoplasm|9814/3|Lymphoma
C569|Ovary|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C569|Ovary|981|Neoplasm|9816/3|Hypodiploid_ALL
C569|Ovary|981|Neoplasm|9817/3|Lymphoma
C569|Ovary|981|Neoplasm|9818/3|Lymphoma
C569|Ovary|981|Neoplasm|9819/3|Leukemia__B_Cell
C569|Ovary|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C569|Ovary|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C569|Ovary|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C569|Ovary|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C569|Ovary|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C569|Ovary|997|Neoplasm|9971/3|Polymorphic_PTLD
C569|Ovary|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C570|Fallopian_Tube|800|Neoplasm|8000/3|Malignant_Neoplasm
C570|Fallopian_Tube|800|Neoplasm|8001/3|Malignant_Cell
C570|Fallopian_Tube|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C570|Fallopian_Tube|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C570|Fallopian_Tube|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C570|Fallopian_Tube|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C570|Fallopian_Tube|801|Carcinoma|8010/2|In_Situ_Cancer
C570|Fallopian_Tube|801|Carcinoma|8010/3|Carcinoma
C570|Fallopian_Tube|801|Carcinoma|8011/3|Malignant_Epithelioma
C570|Fallopian_Tube|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C570|Fallopian_Tube|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C570|Fallopian_Tube|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C570|Fallopian_Tube|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C570|Fallopian_Tube|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C570|Fallopian_Tube|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C570|Fallopian_Tube|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C570|Fallopian_Tube|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C570|Fallopian_Tube|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C570|Fallopian_Tube|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C570|Fallopian_Tube|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C570|Fallopian_Tube|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C570|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C570|Fallopian_Tube|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C570|Fallopian_Tube|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C570|Fallopian_Tube|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C570|Fallopian_Tube|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C570|Fallopian_Tube|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C570|Fallopian_Tube|814|Adenocarcinoma|8140/3|Adenocarcinoma
C570|Fallopian_Tube|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C570|Fallopian_Tube|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C570|Fallopian_Tube|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C570|Fallopian_Tube|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C570|Fallopian_Tube|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C570|Fallopian_Tube|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C570|Fallopian_Tube|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C570|Fallopian_Tube|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C570|Fallopian_Tube|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C570|Fallopian_Tube|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C570|Fallopian_Tube|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C570|Fallopian_Tube|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C570|Fallopian_Tube|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C570|Fallopian_Tube|838|Carcinoma__Endometrioid|8382/3|Carcinoma__Endometrioid
C570|Fallopian_Tube|838|Carcinoma__Endometrioid|8383/3|Carcinoma__Endometrioid
C570|Fallopian_Tube|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C570|Fallopian_Tube|844|Cystadenocarcinoma|8441/2|Serous_Tubal_Intraepithelial_Carcinoma
C570|Fallopian_Tube|844|Cystadenocarcinoma|8441/3|Serous_Cystadenocarcinoma
C570|Fallopian_Tube|846|Papillary_Serous_Cystadenocarcinoma|8460/3|Papillary_Serous_Cystadenocarcinoma
C570|Fallopian_Tube|846|Papillary_Serous_Cystadenocarcinoma|8461/3|Serous_Surface_Papillary_Carcinoma
C570|Fallopian_Tube|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C570|Fallopian_Tube|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C570|Fallopian_Tube|848|Mucinous_Adenocarcinoma|8482/3|Adenocarcinoma__Endocervical_Type
C570|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C570|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C570|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C570|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C570|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C570|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C570|Fallopian_Tube|880|Sarcoma|8800/3|Sarcoma
C570|Fallopian_Tube|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C570|Fallopian_Tube|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C570|Fallopian_Tube|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C570|Fallopian_Tube|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C570|Fallopian_Tube|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C570|Fallopian_Tube|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C570|Fallopian_Tube|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C570|Fallopian_Tube|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C570|Fallopian_Tube|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C570|Fallopian_Tube|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C570|Fallopian_Tube|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C570|Fallopian_Tube|882|Sarcoma|8825/3|Sarcoma
C570|Fallopian_Tube|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C570|Fallopian_Tube|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C570|Fallopian_Tube|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C570|Fallopian_Tube|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C570|Fallopian_Tube|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C570|Fallopian_Tube|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C570|Fallopian_Tube|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C570|Fallopian_Tube|898|Carcinosarcoma|8980/3|Carcinosarcoma
C570|Fallopian_Tube|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C570|Fallopian_Tube|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C570|Fallopian_Tube|911|Mesonephroma|9110/3|Mesonephroma
C570|Fallopian_Tube|959|Lymphoma|9590/3|Lymphoma
C570|Fallopian_Tube|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C570|Fallopian_Tube|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C570|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C570|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C570|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C570|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C570|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C570|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C570|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C570|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C570|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C570|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C570|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C570|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C570|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C570|Fallopian_Tube|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C570|Fallopian_Tube|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C570|Fallopian_Tube|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C570|Fallopian_Tube|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C570|Fallopian_Tube|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C570|Fallopian_Tube|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C570|Fallopian_Tube|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C570|Fallopian_Tube|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C570|Fallopian_Tube|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C570|Fallopian_Tube|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C570|Fallopian_Tube|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C570|Fallopian_Tube|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C570|Fallopian_Tube|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C570|Fallopian_Tube|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C570|Fallopian_Tube|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C570|Fallopian_Tube|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C570|Fallopian_Tube|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C570|Fallopian_Tube|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C570|Fallopian_Tube|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C570|Fallopian_Tube|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C570|Fallopian_Tube|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C570|Fallopian_Tube|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C570|Fallopian_Tube|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C570|Fallopian_Tube|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C570|Fallopian_Tube|973|Plasmacytoma|9731/3|Plasmacytoma
C570|Fallopian_Tube|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C570|Fallopian_Tube|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C570|Fallopian_Tube|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C570|Fallopian_Tube|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C570|Fallopian_Tube|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C570|Fallopian_Tube|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C570|Fallopian_Tube|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C570|Fallopian_Tube|975|Neoplasm|9750/3|Malignant_Histiocytosis
C570|Fallopian_Tube|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C570|Fallopian_Tube|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C570|Fallopian_Tube|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C570|Fallopian_Tube|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C570|Fallopian_Tube|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C570|Fallopian_Tube|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C570|Fallopian_Tube|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C570|Fallopian_Tube|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C570|Fallopian_Tube|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C570|Fallopian_Tube|981|Neoplasm|9812/3|Lymphoma
C570|Fallopian_Tube|981|Neoplasm|9813/3|Lymphoma
C570|Fallopian_Tube|981|Neoplasm|9814/3|Lymphoma
C570|Fallopian_Tube|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C570|Fallopian_Tube|981|Neoplasm|9816/3|Hypodiploid_ALL
C570|Fallopian_Tube|981|Neoplasm|9817/3|Lymphoma
C570|Fallopian_Tube|981|Neoplasm|9818/3|Lymphoma
C570|Fallopian_Tube|981|Neoplasm|9819/3|Leukemia__B_Cell
C570|Fallopian_Tube|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C570|Fallopian_Tube|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C570|Fallopian_Tube|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C570|Fallopian_Tube|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C570|Fallopian_Tube|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C570|Fallopian_Tube|997|Neoplasm|9971/3|Polymorphic_PTLD
C570|Fallopian_Tube|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C571-C574,C577-C579|Fallopian_Tube|800|Neoplasm|8000/3|Malignant_Neoplasm
C571-C574,C577-C579|Fallopian_Tube|800|Neoplasm|8001/3|Malignant_Cell
C571-C574,C577-C579|Fallopian_Tube|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C571-C574,C577-C579|Fallopian_Tube|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C571-C574,C577-C579|Fallopian_Tube|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C571-C574,C577-C579|Fallopian_Tube|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C571-C574,C577-C579|Fallopian_Tube|801|Carcinoma|8010/2|In_Situ_Cancer
C571-C574,C577-C579|Fallopian_Tube|801|Carcinoma|8010/3|Carcinoma
C571-C574,C577-C579|Fallopian_Tube|801|Carcinoma|8011/3|Malignant_Epithelioma
C571-C574,C577-C579|Fallopian_Tube|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C571-C574,C577-C579|Fallopian_Tube|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C571-C574,C577-C579|Fallopian_Tube|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C571-C574,C577-C579|Fallopian_Tube|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C571-C574,C577-C579|Fallopian_Tube|814|Adenocarcinoma|8140/3|Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C571-C574,C577-C579|Fallopian_Tube|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C571-C574,C577-C579|Fallopian_Tube|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C571-C574,C577-C579|Fallopian_Tube|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C571-C574,C577-C579|Fallopian_Tube|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C571-C574,C577-C579|Fallopian_Tube|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C571-C574,C577-C579|Fallopian_Tube|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C571-C574,C577-C579|Fallopian_Tube|838|Carcinoma__Endometrioid|8382/3|Carcinoma__Endometrioid
C571-C574,C577-C579|Fallopian_Tube|838|Carcinoma__Endometrioid|8383/3|Carcinoma__Endometrioid
C571-C574,C577-C579|Fallopian_Tube|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|848|Mucinous_Adenocarcinoma|8482/3|Adenocarcinoma__Endocervical_Type
C571-C574,C577-C579|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C571-C574,C577-C579|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C571-C574,C577-C579|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C571-C574,C577-C579|Fallopian_Tube|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C571-C574,C577-C579|Fallopian_Tube|880|Sarcoma|8800/3|Sarcoma
C571-C574,C577-C579|Fallopian_Tube|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C571-C574,C577-C579|Fallopian_Tube|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C571-C574,C577-C579|Fallopian_Tube|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C571-C574,C577-C579|Fallopian_Tube|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C571-C574,C577-C579|Fallopian_Tube|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C571-C574,C577-C579|Fallopian_Tube|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C571-C574,C577-C579|Fallopian_Tube|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C571-C574,C577-C579|Fallopian_Tube|882|Sarcoma|8825/3|Sarcoma
C571-C574,C577-C579|Fallopian_Tube|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C571-C574,C577-C579|Fallopian_Tube|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C571-C574,C577-C579|Fallopian_Tube|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C571-C574,C577-C579|Fallopian_Tube|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C571-C574,C577-C579|Fallopian_Tube|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C571-C574,C577-C579|Fallopian_Tube|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C571-C574,C577-C579|Fallopian_Tube|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C571-C574,C577-C579|Fallopian_Tube|898|Carcinosarcoma|8980/3|Carcinosarcoma
C571-C574,C577-C579|Fallopian_Tube|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C571-C574,C577-C579|Fallopian_Tube|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C571-C574,C577-C579|Fallopian_Tube|911|Mesonephroma|9110/3|Mesonephroma
C571-C574,C577-C579|Fallopian_Tube|959|Lymphoma|9590/3|Lymphoma
C571-C574,C577-C579|Fallopian_Tube|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C571-C574,C577-C579|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C571-C574,C577-C579|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C571-C574,C577-C579|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C571-C574,C577-C579|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C571-C574,C577-C579|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C571-C574,C577-C579|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C571-C574,C577-C579|Fallopian_Tube|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C571-C574,C577-C579|Fallopian_Tube|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C571-C574,C577-C579|Fallopian_Tube|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C571-C574,C577-C579|Fallopian_Tube|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C571-C574,C577-C579|Fallopian_Tube|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C571-C574,C577-C579|Fallopian_Tube|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C571-C574,C577-C579|Fallopian_Tube|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|973|Plasmacytoma|9731/3|Plasmacytoma
C571-C574,C577-C579|Fallopian_Tube|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C571-C574,C577-C579|Fallopian_Tube|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C571-C574,C577-C579|Fallopian_Tube|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C571-C574,C577-C579|Fallopian_Tube|975|Neoplasm|9750/3|Malignant_Histiocytosis
C571-C574,C577-C579|Fallopian_Tube|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C571-C574,C577-C579|Fallopian_Tube|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C571-C574,C577-C579|Fallopian_Tube|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C571-C574,C577-C579|Fallopian_Tube|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C571-C574,C577-C579|Fallopian_Tube|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9812/3|Lymphoma
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9813/3|Lymphoma
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9814/3|Lymphoma
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9816/3|Hypodiploid_ALL
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9817/3|Lymphoma
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9818/3|Lymphoma
C571-C574,C577-C579|Fallopian_Tube|981|Neoplasm|9819/3|Leukemia__B_Cell
C571-C574,C577-C579|Fallopian_Tube|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C571-C574,C577-C579|Fallopian_Tube|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C571-C574,C577-C579|Fallopian_Tube|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C571-C574,C577-C579|Fallopian_Tube|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C571-C574,C577-C579|Fallopian_Tube|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C571-C574,C577-C579|Fallopian_Tube|997|Neoplasm|9971/3|Polymorphic_PTLD
C571-C574,C577-C579|Fallopian_Tube|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C589|Placenta_Part|800|Neoplasm|8000/3|Malignant_Neoplasm
C589|Placenta_Part|800|Neoplasm|8001/3|Malignant_Cell
C589|Placenta_Part|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C589|Placenta_Part|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C589|Placenta_Part|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C589|Placenta_Part|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C589|Placenta_Part|910|Choriocarcinoma|9100/3|Choriocarcinoma
C589|Placenta_Part|910|Choriocarcinoma|9101/3|Choriocarcinoma
C589|Placenta_Part|910|Choriocarcinoma|9104/3|Placental_Site_GTT
C589|Placenta_Part|910|Choriocarcinoma|9105/3|Epithelioid_Trophoblastic_Tumor
C589|Placenta_Part|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C589|Placenta_Part|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C600-C602,C608-C609|Penis|800|Neoplasm|8000/3|Malignant_Neoplasm
C600-C602,C608-C609|Penis|800|Neoplasm|8001/3|Malignant_Cell
C600-C602,C608-C609|Penis|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C600-C602,C608-C609|Penis|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C600-C602,C608-C609|Penis|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C600-C602,C608-C609|Penis|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C600-C602,C608-C609|Penis|801|Carcinoma|8010/2|In_Situ_Cancer
C600-C602,C608-C609|Penis|801|Carcinoma|8010/3|Carcinoma
C600-C602,C608-C609|Penis|801|Carcinoma|8011/3|Malignant_Epithelioma
C600-C602,C608-C609|Penis|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C600-C602,C608-C609|Penis|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C600-C602,C608-C609|Penis|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C600-C602,C608-C609|Penis|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C600-C602,C608-C609|Penis|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C600-C602,C608-C609|Penis|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C600-C602,C608-C609|Penis|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C600-C602,C608-C609|Penis|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C600-C602,C608-C609|Penis|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C600-C602,C608-C609|Penis|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C600-C602,C608-C609|Penis|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|805|Papillary_Carcinoma|8054/3|Verrucous_Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8071/2|Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C600-C602,C608-C609|Penis|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|808|Lymphoepithelial_Carcinoma|8080/2|Penile_Carcinoma_In_Situ
C600-C602,C608-C609|Penis|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C600-C602,C608-C609|Penis|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C600-C602,C608-C609|Penis|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|809|Basal_Cell_Carcinoma|8090/3|Basal_Cell_Carcinoma
C600-C602,C608-C609|Penis|809|Basal_Cell_Carcinoma|8091/3|Superficial_Basal_Cell_Carcinoma
C600-C602,C608-C609|Penis|809|Basal_Cell_Carcinoma|8092/3|Skin_Infiltrating_Basal_Cell_Carcinoma
C600-C602,C608-C609|Penis|809|Basal_Cell_Carcinoma|8093/3|Fibroepithelioma_Of_Pinkus
C600-C602,C608-C609|Penis|809|Basal_Cell_Carcinoma|8094/3|Skin_Basosquamous_Cell_Carcinoma
C600-C602,C608-C609|Penis|809|Basal_Cell_Carcinoma|8095/3|Skin_Metatypical_Carcinoma
C600-C602,C608-C609|Penis|809|Basal_Cell_Carcinoma|8097/3|Skin_Nodular_Basal_Cell_Carcinoma
C600-C602,C608-C609|Penis|809|Basal_Cell_Carcinoma|8098/3|Skin_Adenoid_Basal_Cell_Carcinoma
C600-C602,C608-C609|Penis|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C600-C602,C608-C609|Penis|811|Pilomatrical_Carcinoma|8110/3|Pilomatrical_Carcinoma
C600-C602,C608-C609|Penis|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C600-C602,C608-C609|Penis|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C600-C602,C608-C609|Penis|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C600-C602,C608-C609|Penis|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C600-C602,C608-C609|Penis|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C600-C602,C608-C609|Penis|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8140/3|Adenocarcinoma
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C600-C602,C608-C609|Penis|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C600-C602,C608-C609|Penis|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C600-C602,C608-C609|Penis|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C600-C602,C608-C609|Penis|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C600-C602,C608-C609|Penis|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C600-C602,C608-C609|Penis|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C600-C602,C608-C609|Penis|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C600-C602,C608-C609|Penis|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C600-C602,C608-C609|Penis|839|Adnexal_Carcinoma|8390/3|Adnexal_Carcinoma
C600-C602,C608-C609|Penis|840|Sweat_Gland_Adenocarcinoma|8400/3|Sweat_Gland_Adenocarcinoma
C600-C602,C608-C609|Penis|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C600-C602,C608-C609|Penis|841|Eccrine_Adenocarcinoma|8410/3|Sebaceous_Adenocarcinoma
C600-C602,C608-C609|Penis|841|Eccrine_Adenocarcinoma|8413/3|Eccrine_Adenocarcinoma
C600-C602,C608-C609|Penis|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C600-C602,C608-C609|Penis|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C600-C602,C608-C609|Penis|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C600-C602,C608-C609|Penis|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C600-C602,C608-C609|Penis|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C600-C602,C608-C609|Penis|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C600-C602,C608-C609|Penis|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C600-C602,C608-C609|Penis|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C600-C602,C608-C609|Penis|872|Melanoma|8720/3|Melanoma
C600-C602,C608-C609|Penis|872|Melanoma|8721/3|Nodular_Melanoma
C600-C602,C608-C609|Penis|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C600-C602,C608-C609|Penis|872|Melanoma|8723/3|Regressing_Melanoma
C600-C602,C608-C609|Penis|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C600-C602,C608-C609|Penis|874|Nevus|8740/3|Melanoma_In_Junctional_Nevus
C600-C602,C608-C609|Penis|874|Nevus|8741/2|Precancerous_Melanosis
C600-C602,C608-C609|Penis|874|Nevus|8741/3|Melanoma
C600-C602,C608-C609|Penis|874|Nevus|8742/2|Lentigo_Maligna
C600-C602,C608-C609|Penis|874|Nevus|8742/3|Lentigo_Maligna_Melanoma
C600-C602,C608-C609|Penis|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C600-C602,C608-C609|Penis|874|Nevus|8745/3|Desmoplastic_Melanoma
C600-C602,C608-C609|Penis|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C600-C602,C608-C609|Penis|876|Nevus|8761/3|Giant_Congenital_Nevus
C600-C602,C608-C609|Penis|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C600-C602,C608-C609|Penis|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C600-C602,C608-C609|Penis|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C600-C602,C608-C609|Penis|878|Melanoma_Arising_From_Blue_Nevus|8780/3|Melanoma_Arising_From_Blue_Nevus
C600-C602,C608-C609|Penis|880|Sarcoma|8800/3|Sarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C600-C602,C608-C609|Penis|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C600-C602,C608-C609|Penis|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C600-C602,C608-C609|Penis|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C600-C602,C608-C609|Penis|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C600-C602,C608-C609|Penis|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C600-C602,C608-C609|Penis|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C600-C602,C608-C609|Penis|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C600-C602,C608-C609|Penis|882|Sarcoma|8825/3|Sarcoma
C600-C602,C608-C609|Penis|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8850/3|Liposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C600-C602,C608-C609|Penis|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8855/3|Liposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C600-C602,C608-C609|Penis|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C600-C602,C608-C609|Penis|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C600-C602,C608-C609|Penis|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C600-C602,C608-C609|Penis|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C600-C602,C608-C609|Penis|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C600-C602,C608-C609|Penis|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C600-C602,C608-C609|Penis|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C600-C602,C608-C609|Penis|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C600-C602,C608-C609|Penis|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C600-C602,C608-C609|Penis|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C600-C602,C608-C609|Penis|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C600-C602,C608-C609|Penis|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C600-C602,C608-C609|Penis|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C600-C602,C608-C609|Penis|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C600-C602,C608-C609|Penis|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C600-C602,C608-C609|Penis|898|Carcinosarcoma|8980/3|Carcinosarcoma
C600-C602,C608-C609|Penis|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C600-C602,C608-C609|Penis|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C600-C602,C608-C609|Penis|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C600-C602,C608-C609|Penis|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C600-C602,C608-C609|Penis|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C600-C602,C608-C609|Penis|959|Lymphoma|9597/3|Crosti_s_Disease
C600-C602,C608-C609|Penis|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C600-C602,C608-C609|Penis|970|T_Cell_Lymphoma|9700/3|Mycosis_Fungoides
C600-C602,C608-C609|Penis|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C600-C602,C608-C609|Penis|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C600-C602,C608-C609|Penis|970|T_Cell_Lymphoma|9709/3|Cutaneous_T_Cell_Non_Hodgkin_Lymphoma
C600-C602,C608-C609|Penis|971|Adult_Non_Hodgkin_Lymphoma|9718/3|C_ALCL
C600-C602,C608-C609|Penis|972|Lymphoblastic_Lymphoma|9725/3|Hydroa_Vacciniforme_Like_Lymphoma
C600-C602,C608-C609|Penis|972|Lymphoblastic_Lymphoma|9726/3|T_Cell_Lymphoma
C600-C602,C608-C609|Penis|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C619|Prostate|800|Neoplasm|8000/3|Malignant_Neoplasm
C619|Prostate|800|Neoplasm|8001/3|Malignant_Cell
C619|Prostate|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C619|Prostate|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C619|Prostate|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C619|Prostate|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C619|Prostate|801|Carcinoma|8010/2|In_Situ_Cancer
C619|Prostate|801|Carcinoma|8010/3|Carcinoma
C619|Prostate|801|Carcinoma|8011/3|Malignant_Epithelioma
C619|Prostate|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C619|Prostate|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C619|Prostate|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C619|Prostate|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C619|Prostate|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C619|Prostate|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C619|Prostate|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C619|Prostate|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C619|Prostate|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C619|Prostate|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C619|Prostate|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C619|Prostate|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C619|Prostate|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C619|Prostate|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C619|Prostate|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C619|Prostate|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C619|Prostate|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C619|Prostate|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C619|Prostate|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C619|Prostate|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C619|Prostate|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C619|Prostate|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C619|Prostate|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C619|Prostate|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C619|Prostate|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C619|Prostate|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C619|Prostate|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C619|Prostate|813|Carcinoma|8130/2|Carcinoma
C619|Prostate|813|Carcinoma|8130/3|Carcinoma
C619|Prostate|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C619|Prostate|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C619|Prostate|814|Adenocarcinoma|8140/3|Adenocarcinoma
C619|Prostate|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C619|Prostate|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C619|Prostate|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C619|Prostate|814|Adenocarcinoma|8148/2|Intraepithelial_Neoplasia
C619|Prostate|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C619|Prostate|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C619|Prostate|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C619|Prostate|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C619|Prostate|825|Bronchioloalveolar_Adenocarcinoma|8251/3|Bronchioloalveolar_Adenocarcinoma
C619|Prostate|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C619|Prostate|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C619|Prostate|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C619|Prostate|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C619|Prostate|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C619|Prostate|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C619|Prostate|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C619|Prostate|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C619|Prostate|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C619|Prostate|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C619|Prostate|850|Ductal_Carcinoma|8500/2|Ductal_Breast_Carcinoma_In_Situ
C619|Prostate|850|Ductal_Carcinoma|8500/3|Invasive_Carcinoma
C619|Prostate|850|Ductal_Carcinoma|8503/2|Intraductal_Papillary_Breast_Carcinoma
C619|Prostate|850|Ductal_Carcinoma|8503/3|Intraductal_Papillary_Breast_Carcinoma
C619|Prostate|850|Ductal_Carcinoma|8504/2|Intracystic_Papillary_Breast_Carcinoma
C619|Prostate|850|Ductal_Carcinoma|8504/3|Intracystic_Papillary_Breast_Carcinoma
C619|Prostate|850|Ductal_Carcinoma|8507/2|Micropapillary_Carcinoma
C619|Prostate|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C619|Prostate|851|Medullary_Carcinoma|8514/3|Ductal_Carcinoma
C619|Prostate|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C619|Prostate|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C619|Prostate|855|Acinar_Cell_Carcinoma|8552/3|Ductal_Carcinoma
C619|Prostate|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C619|Prostate|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C619|Prostate|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C619|Prostate|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C619|Prostate|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C619|Prostate|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C619|Prostate|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C619|Prostate|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C619|Prostate|880|Sarcoma|8800/3|Sarcoma
C619|Prostate|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C619|Prostate|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C619|Prostate|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C619|Prostate|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C619|Prostate|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C619|Prostate|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C619|Prostate|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C619|Prostate|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C619|Prostate|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C619|Prostate|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C619|Prostate|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C619|Prostate|882|Sarcoma|8825/3|Sarcoma
C619|Prostate|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C619|Prostate|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C619|Prostate|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C619|Prostate|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C619|Prostate|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C619|Prostate|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C619|Prostate|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C619|Prostate|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C619|Prostate|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C619|Prostate|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C619|Prostate|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C619|Prostate|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C619|Prostate|898|Carcinosarcoma|8980/3|Carcinosarcoma
C619|Prostate|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C619|Prostate|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C619|Prostate|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C619|Prostate|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C619|Prostate|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C619|Prostate|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C619|Prostate|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C619|Prostate|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C619|Prostate|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C619|Prostate|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C619|Prostate|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C619|Prostate|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C619|Prostate|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C619|Prostate|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C619|Prostate|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C619|Prostate|981|Neoplasm|9812/3|Lymphoma
C619|Prostate|981|Neoplasm|9813/3|Lymphoma
C619|Prostate|981|Neoplasm|9814/3|Lymphoma
C619|Prostate|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C619|Prostate|981|Neoplasm|9816/3|Hypodiploid_ALL
C619|Prostate|981|Neoplasm|9817/3|Lymphoma
C619|Prostate|981|Neoplasm|9818/3|Lymphoma
C619|Prostate|981|Neoplasm|9819/3|Leukemia__B_Cell
C619|Prostate|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C619|Prostate|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C619|Prostate|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C619|Prostate|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C619|Prostate|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C619|Prostate|997|Neoplasm|9971/3|Polymorphic_PTLD
C619|Prostate|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C620-C621,C629|Testis|800|Neoplasm|8000/3|Malignant_Neoplasm
C620-C621,C629|Testis|800|Neoplasm|8001/3|Malignant_Cell
C620-C621,C629|Testis|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C620-C621,C629|Testis|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C620-C621,C629|Testis|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C620-C621,C629|Testis|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C620-C621,C629|Testis|801|Carcinoma|8010/2|In_Situ_Cancer
C620-C621,C629|Testis|801|Carcinoma|8010/3|Carcinoma
C620-C621,C629|Testis|801|Carcinoma|8011/3|Malignant_Epithelioma
C620-C621,C629|Testis|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C620-C621,C629|Testis|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C620-C621,C629|Testis|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C620-C621,C629|Testis|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C620-C621,C629|Testis|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C620-C621,C629|Testis|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C620-C621,C629|Testis|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C620-C621,C629|Testis|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C620-C621,C629|Testis|814|Adenocarcinoma|8140/3|Adenocarcinoma
C620-C621,C629|Testis|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C620-C621,C629|Testis|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C620-C621,C629|Testis|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C620-C621,C629|Testis|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C620-C621,C629|Testis|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C620-C621,C629|Testis|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C620-C621,C629|Testis|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C620-C621,C629|Testis|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C620-C621,C629|Testis|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C620-C621,C629|Testis|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C620-C621,C629|Testis|863|Neoplasm|8630/3|Malignant_Sertoli_Cell_Tumor
C620-C621,C629|Testis|863|Neoplasm|8631/3|Sertoli_Leydig_Cell_Tumor
C620-C621,C629|Testis|863|Neoplasm|8634/3|Sertoli_Leydig_Cell_Tumor
C620-C621,C629|Testis|864|Sertoli_Cell_Carcinoma|8640/3|Sertoli_Cell_Carcinoma
C620-C621,C629|Testis|865|Malignant_Leydig_Cell_Tumor|8650/3|Malignant_Leydig_Cell_Tumor
C620-C621,C629|Testis|880|Sarcoma|8800/3|Sarcoma
C620-C621,C629|Testis|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C620-C621,C629|Testis|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C620-C621,C629|Testis|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C620-C621,C629|Testis|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C620-C621,C629|Testis|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C620-C621,C629|Testis|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C620-C621,C629|Testis|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C620-C621,C629|Testis|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C620-C621,C629|Testis|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C620-C621,C629|Testis|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C620-C621,C629|Testis|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C620-C621,C629|Testis|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C620-C621,C629|Testis|906|Germ_Cell_Tumor|9061/3|Seminoma
C620-C621,C629|Testis|906|Germ_Cell_Tumor|9062/3|Atypical_Seminoma
C620-C621,C629|Testis|906|Germ_Cell_Tumor|9063/3|Testicular_Spermatocytic_Seminoma
C620-C621,C629|Testis|906|Germ_Cell_Tumor|9064/2|Intratubular_Germ_Cell_Neoplasia
C620-C621,C629|Testis|906|Germ_Cell_Tumor|9064/3|Germinoma
C620-C621,C629|Testis|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C620-C621,C629|Testis|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C620-C621,C629|Testis|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C620-C621,C629|Testis|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C620-C621,C629|Testis|908|Teratoma|9080/3|Immature_Teratoma
C620-C621,C629|Testis|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C620-C621,C629|Testis|908|Teratoma|9082/3|Immature_Teratoma
C620-C621,C629|Testis|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C620-C621,C629|Testis|908|Teratoma|9084/3|Teratoma
C620-C621,C629|Testis|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C620-C621,C629|Testis|910|Choriocarcinoma|9100/3|Choriocarcinoma
C620-C621,C629|Testis|910|Choriocarcinoma|9101/3|Choriocarcinoma
C620-C621,C629|Testis|910|Choriocarcinoma|9102/3|Malignant_Trophoblastic_Teratoma
C620-C621,C629|Testis|910|Choriocarcinoma|9105/3|Epithelioid_Trophoblastic_Tumor
C620-C621,C629|Testis|959|Lymphoma|9590/3|Lymphoma
C620-C621,C629|Testis|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C620-C621,C629|Testis|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C620-C621,C629|Testis|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C620-C621,C629|Testis|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C620-C621,C629|Testis|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C620-C621,C629|Testis|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C620-C621,C629|Testis|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C620-C621,C629|Testis|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C620-C621,C629|Testis|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C620-C621,C629|Testis|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C620-C621,C629|Testis|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C620-C621,C629|Testis|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C620-C621,C629|Testis|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C620-C621,C629|Testis|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C620-C621,C629|Testis|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C620-C621,C629|Testis|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C620-C621,C629|Testis|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C620-C621,C629|Testis|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C620-C621,C629|Testis|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C620-C621,C629|Testis|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C620-C621,C629|Testis|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C620-C621,C629|Testis|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C620-C621,C629|Testis|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C620-C621,C629|Testis|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C620-C621,C629|Testis|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C620-C621,C629|Testis|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C620-C621,C629|Testis|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C620-C621,C629|Testis|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C620-C621,C629|Testis|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C620-C621,C629|Testis|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C620-C621,C629|Testis|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C620-C621,C629|Testis|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C620-C621,C629|Testis|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C620-C621,C629|Testis|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C620-C621,C629|Testis|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C620-C621,C629|Testis|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C620-C621,C629|Testis|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C620-C621,C629|Testis|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C620-C621,C629|Testis|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C620-C621,C629|Testis|973|Plasmacytoma|9731/3|Plasmacytoma
C620-C621,C629|Testis|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C620-C621,C629|Testis|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C620-C621,C629|Testis|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C620-C621,C629|Testis|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C620-C621,C629|Testis|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C620-C621,C629|Testis|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C620-C621,C629|Testis|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C620-C621,C629|Testis|975|Neoplasm|9750/3|Malignant_Histiocytosis
C620-C621,C629|Testis|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C620-C621,C629|Testis|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C620-C621,C629|Testis|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C620-C621,C629|Testis|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C620-C621,C629|Testis|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C620-C621,C629|Testis|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C620-C621,C629|Testis|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C620-C621,C629|Testis|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C620-C621,C629|Testis|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C620-C621,C629|Testis|981|Neoplasm|9812/3|Lymphoma
C620-C621,C629|Testis|981|Neoplasm|9813/3|Lymphoma
C620-C621,C629|Testis|981|Neoplasm|9814/3|Lymphoma
C620-C621,C629|Testis|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C620-C621,C629|Testis|981|Neoplasm|9816/3|Hypodiploid_ALL
C620-C621,C629|Testis|981|Neoplasm|9817/3|Lymphoma
C620-C621,C629|Testis|981|Neoplasm|9818/3|Lymphoma
C620-C621,C629|Testis|981|Neoplasm|9819/3|Leukemia__B_Cell
C620-C621,C629|Testis|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C620-C621,C629|Testis|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C620-C621,C629|Testis|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C620-C621,C629|Testis|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C620-C621,C629|Testis|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C620-C621,C629|Testis|997|Neoplasm|9971/3|Polymorphic_PTLD
C620-C621,C629|Testis|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C630, C631, C637-C639|Spermatic_Cord|800|Neoplasm|8000/3|Malignant_Neoplasm
C630, C631, C637-C639|Spermatic_Cord|800|Neoplasm|8001/3|Malignant_Cell
C630, C631, C637-C639|Spermatic_Cord|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C630, C631, C637-C639|Spermatic_Cord|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C630, C631, C637-C639|Spermatic_Cord|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C630, C631, C637-C639|Spermatic_Cord|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C630, C631, C637-C639|Spermatic_Cord|801|Carcinoma|8010/2|In_Situ_Cancer
C630, C631, C637-C639|Spermatic_Cord|801|Carcinoma|8010/3|Carcinoma
C630, C631, C637-C639|Spermatic_Cord|801|Carcinoma|8011/3|Malignant_Epithelioma
C630, C631, C637-C639|Spermatic_Cord|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C630, C631, C637-C639|Spermatic_Cord|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C630, C631, C637-C639|Spermatic_Cord|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C630, C631, C637-C639|Spermatic_Cord|814|Adenocarcinoma|8140/3|Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C630, C631, C637-C639|Spermatic_Cord|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C630, C631, C637-C639|Spermatic_Cord|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C630, C631, C637-C639|Spermatic_Cord|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C630, C631, C637-C639|Spermatic_Cord|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C630, C631, C637-C639|Spermatic_Cord|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C630, C631, C637-C639|Spermatic_Cord|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C630, C631, C637-C639|Spermatic_Cord|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C630, C631, C637-C639|Spermatic_Cord|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C630, C631, C637-C639|Spermatic_Cord|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C630, C631, C637-C639|Spermatic_Cord|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C630, C631, C637-C639|Spermatic_Cord|880|Sarcoma|8800/3|Sarcoma
C630, C631, C637-C639|Spermatic_Cord|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C630, C631, C637-C639|Spermatic_Cord|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C630, C631, C637-C639|Spermatic_Cord|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C630, C631, C637-C639|Spermatic_Cord|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C630, C631, C637-C639|Spermatic_Cord|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C630, C631, C637-C639|Spermatic_Cord|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C630, C631, C637-C639|Spermatic_Cord|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C630, C631, C637-C639|Spermatic_Cord|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C630, C631, C637-C639|Spermatic_Cord|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C630, C631, C637-C639|Spermatic_Cord|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C630, C631, C637-C639|Spermatic_Cord|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C630, C631, C637-C639|Spermatic_Cord|882|Sarcoma|8825/3|Sarcoma
C630, C631, C637-C639|Spermatic_Cord|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C630, C631, C637-C639|Spermatic_Cord|885|Liposarcoma|8850/3|Liposarcoma
C630, C631, C637-C639|Spermatic_Cord|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C630, C631, C637-C639|Spermatic_Cord|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C630, C631, C637-C639|Spermatic_Cord|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C630, C631, C637-C639|Spermatic_Cord|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C630, C631, C637-C639|Spermatic_Cord|885|Liposarcoma|8855/3|Liposarcoma
C630, C631, C637-C639|Spermatic_Cord|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C630, C631, C637-C639|Spermatic_Cord|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C630, C631, C637-C639|Spermatic_Cord|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C630, C631, C637-C639|Spermatic_Cord|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C630, C631, C637-C639|Spermatic_Cord|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C630, C631, C637-C639|Spermatic_Cord|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C630, C631, C637-C639|Spermatic_Cord|898|Carcinosarcoma|8980/3|Carcinosarcoma
C630, C631, C637-C639|Spermatic_Cord|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C630, C631, C637-C639|Spermatic_Cord|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C630, C631, C637-C639|Spermatic_Cord|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C630, C631, C637-C639|Spermatic_Cord|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C630, C631, C637-C639|Spermatic_Cord|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C630, C631, C637-C639|Spermatic_Cord|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C630, C631, C637-C639|Spermatic_Cord|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C632|Scrotum|800|Neoplasm|8000/3|Malignant_Neoplasm
C632|Scrotum|800|Neoplasm|8001/3|Malignant_Cell
C632|Scrotum|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C632|Scrotum|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C632|Scrotum|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C632|Scrotum|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C632|Scrotum|801|Carcinoma|8010/2|In_Situ_Cancer
C632|Scrotum|801|Carcinoma|8010/3|Carcinoma
C632|Scrotum|801|Carcinoma|8011/3|Malignant_Epithelioma
C632|Scrotum|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C632|Scrotum|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C632|Scrotum|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C632|Scrotum|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C632|Scrotum|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C632|Scrotum|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C632|Scrotum|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C632|Scrotum|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C632|Scrotum|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C632|Scrotum|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C632|Scrotum|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C632|Scrotum|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C632|Scrotum|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C632|Scrotum|808|Lymphoepithelial_Carcinoma|8080/2|Penile_Carcinoma_In_Situ
C632|Scrotum|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C632|Scrotum|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C632|Scrotum|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C632|Scrotum|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C632|Scrotum|809|Basal_Cell_Carcinoma|8090/3|Basal_Cell_Carcinoma
C632|Scrotum|809|Basal_Cell_Carcinoma|8091/3|Superficial_Basal_Cell_Carcinoma
C632|Scrotum|809|Basal_Cell_Carcinoma|8092/3|Skin_Infiltrating_Basal_Cell_Carcinoma
C632|Scrotum|809|Basal_Cell_Carcinoma|8093/3|Fibroepithelioma_Of_Pinkus
C632|Scrotum|809|Basal_Cell_Carcinoma|8094/3|Skin_Basosquamous_Cell_Carcinoma
C632|Scrotum|809|Basal_Cell_Carcinoma|8095/3|Skin_Metatypical_Carcinoma
C632|Scrotum|809|Basal_Cell_Carcinoma|8097/3|Skin_Nodular_Basal_Cell_Carcinoma
C632|Scrotum|809|Basal_Cell_Carcinoma|8098/3|Skin_Adenoid_Basal_Cell_Carcinoma
C632|Scrotum|810|Trichilemmocarcinoma|8102/3|Trichilemmocarcinoma
C632|Scrotum|811|Pilomatrical_Carcinoma|8110/3|Pilomatrical_Carcinoma
C632|Scrotum|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C632|Scrotum|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C632|Scrotum|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C632|Scrotum|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C632|Scrotum|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C632|Scrotum|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C632|Scrotum|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C632|Scrotum|814|Adenocarcinoma|8140/3|Adenocarcinoma
C632|Scrotum|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C632|Scrotum|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C632|Scrotum|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C632|Scrotum|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C632|Scrotum|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C632|Scrotum|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C632|Scrotum|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C632|Scrotum|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C632|Scrotum|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C632|Scrotum|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C632|Scrotum|839|Adnexal_Carcinoma|8390/3|Adnexal_Carcinoma
C632|Scrotum|840|Sweat_Gland_Adenocarcinoma|8400/3|Sweat_Gland_Adenocarcinoma
C632|Scrotum|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C632|Scrotum|841|Eccrine_Adenocarcinoma|8410/3|Sebaceous_Adenocarcinoma
C632|Scrotum|841|Eccrine_Adenocarcinoma|8413/3|Eccrine_Adenocarcinoma
C632|Scrotum|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C632|Scrotum|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C632|Scrotum|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C632|Scrotum|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C632|Scrotum|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C632|Scrotum|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C632|Scrotum|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C632|Scrotum|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C632|Scrotum|872|Melanoma|8720/3|Melanoma
C632|Scrotum|872|Melanoma|8721/3|Nodular_Melanoma
C632|Scrotum|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C632|Scrotum|872|Melanoma|8723/3|Regressing_Melanoma
C632|Scrotum|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C632|Scrotum|874|Nevus|8740/3|Melanoma_In_Junctional_Nevus
C632|Scrotum|874|Nevus|8741/2|Precancerous_Melanosis
C632|Scrotum|874|Nevus|8741/3|Melanoma
C632|Scrotum|874|Nevus|8742/2|Lentigo_Maligna
C632|Scrotum|874|Nevus|8742/3|Lentigo_Maligna_Melanoma
C632|Scrotum|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C632|Scrotum|874|Nevus|8745/3|Desmoplastic_Melanoma
C632|Scrotum|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C632|Scrotum|876|Nevus|8761/3|Giant_Congenital_Nevus
C632|Scrotum|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C632|Scrotum|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C632|Scrotum|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C632|Scrotum|878|Melanoma_Arising_From_Blue_Nevus|8780/3|Melanoma_Arising_From_Blue_Nevus
C632|Scrotum|880|Sarcoma|8800/3|Sarcoma
C632|Scrotum|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C632|Scrotum|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C632|Scrotum|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C632|Scrotum|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C632|Scrotum|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C632|Scrotum|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C632|Scrotum|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C632|Scrotum|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C632|Scrotum|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C632|Scrotum|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C632|Scrotum|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C632|Scrotum|882|Sarcoma|8825/3|Sarcoma
C632|Scrotum|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C632|Scrotum|885|Liposarcoma|8850/3|Liposarcoma
C632|Scrotum|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C632|Scrotum|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C632|Scrotum|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C632|Scrotum|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C632|Scrotum|885|Liposarcoma|8855/3|Liposarcoma
C632|Scrotum|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C632|Scrotum|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C632|Scrotum|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C632|Scrotum|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C632|Scrotum|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C632|Scrotum|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C632|Scrotum|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C632|Scrotum|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C632|Scrotum|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C632|Scrotum|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C632|Scrotum|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C632|Scrotum|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C632|Scrotum|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C632|Scrotum|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C632|Scrotum|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C632|Scrotum|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C632|Scrotum|898|Carcinosarcoma|8980/3|Carcinosarcoma
C632|Scrotum|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C632|Scrotum|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C632|Scrotum|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C632|Scrotum|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C632|Scrotum|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C632|Scrotum|959|Lymphoma|9597/3|Crosti_s_Disease
C632|Scrotum|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C632|Scrotum|970|T_Cell_Lymphoma|9700/3|Mycosis_Fungoides
C632|Scrotum|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C632|Scrotum|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C632|Scrotum|970|T_Cell_Lymphoma|9709/3|Cutaneous_T_Cell_Non_Hodgkin_Lymphoma
C632|Scrotum|971|Adult_Non_Hodgkin_Lymphoma|9718/3|C_ALCL
C632|Scrotum|972|Lymphoblastic_Lymphoma|9725/3|Hydroa_Vacciniforme_Like_Lymphoma
C632|Scrotum|972|Lymphoblastic_Lymphoma|9726/3|T_Cell_Lymphoma
C632|Scrotum|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C649|Kidney|800|Neoplasm|8000/3|Malignant_Neoplasm
C649|Kidney|800|Neoplasm|8001/3|Malignant_Cell
C649|Kidney|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C649|Kidney|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C649|Kidney|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C649|Kidney|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C649|Kidney|801|Carcinoma|8010/2|In_Situ_Cancer
C649|Kidney|801|Carcinoma|8010/3|Carcinoma
C649|Kidney|801|Carcinoma|8011/3|Malignant_Epithelioma
C649|Kidney|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C649|Kidney|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C649|Kidney|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C649|Kidney|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C649|Kidney|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C649|Kidney|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C649|Kidney|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C649|Kidney|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C649|Kidney|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C649|Kidney|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C649|Kidney|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C649|Kidney|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C649|Kidney|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C649|Kidney|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C649|Kidney|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C649|Kidney|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C649|Kidney|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C649|Kidney|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C649|Kidney|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C649|Kidney|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C649|Kidney|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C649|Kidney|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C649|Kidney|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C649|Kidney|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C649|Kidney|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C649|Kidney|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C649|Kidney|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C649|Kidney|813|Carcinoma|8130/2|Carcinoma
C649|Kidney|813|Carcinoma|8130/3|Carcinoma
C649|Kidney|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C649|Kidney|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C649|Kidney|814|Adenocarcinoma|8140/3|Adenocarcinoma
C649|Kidney|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C649|Kidney|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C649|Kidney|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C649|Kidney|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C649|Kidney|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C649|Kidney|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C649|Kidney|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C649|Kidney|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C649|Kidney|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C649|Kidney|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C649|Kidney|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C649|Kidney|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C649|Kidney|831|Clear_Cell_Adenocarcinoma|8311/3|Renal_Cell_Carcinoma
C649|Kidney|831|Clear_Cell_Adenocarcinoma|8312/3|Renal_Cell_Carcinoma
C649|Kidney|831|Clear_Cell_Adenocarcinoma|8316/3|Cyst_associated_Renal_Cell_Carcinoma
C649|Kidney|831|Clear_Cell_Adenocarcinoma|8317/3|Chromophobe_Renal_Cell_Carcinoma
C649|Kidney|831|Clear_Cell_Adenocarcinoma|8318/3|Sarcomatoid_Renal_Cell_Carcinoma
C649|Kidney|831|Clear_Cell_Adenocarcinoma|8319/3|Collecting_Duct_Carcinoma_Of_Kidney
C649|Kidney|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C649|Kidney|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C649|Kidney|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C649|Kidney|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C649|Kidney|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C649|Kidney|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C649|Kidney|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C649|Kidney|880|Sarcoma|8800/3|Sarcoma
C649|Kidney|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C649|Kidney|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C649|Kidney|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C649|Kidney|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C649|Kidney|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C649|Kidney|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C649|Kidney|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C649|Kidney|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C649|Kidney|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C649|Kidney|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C649|Kidney|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C649|Kidney|882|Sarcoma|8825/3|Sarcoma
C649|Kidney|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C649|Kidney|885|Liposarcoma|8850/3|Liposarcoma
C649|Kidney|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C649|Kidney|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C649|Kidney|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C649|Kidney|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C649|Kidney|885|Liposarcoma|8855/3|Liposarcoma
C649|Kidney|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C649|Kidney|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C649|Kidney|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C649|Kidney|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C649|Kidney|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C649|Kidney|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C649|Kidney|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C649|Kidney|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C649|Kidney|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C649|Kidney|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C649|Kidney|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C649|Kidney|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C649|Kidney|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C649|Kidney|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C649|Kidney|895|Mixed_Tumor__Mullerian|8959/3|Malignant_Cystic_Nephroma
C649|Kidney|896|Nephroblastoma|8960/3|Nephroblastoma
C649|Kidney|896|Nephroblastoma|8963/3|Rhabdoid_Tumor
C649|Kidney|896|Nephroblastoma|8964/3|Clear_Cell_Sarcoma_Of_The_Kidney
C649|Kidney|898|Carcinosarcoma|8980/3|Carcinosarcoma
C649|Kidney|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C649|Kidney|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C649|Kidney|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C649|Kidney|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C649|Kidney|950|Neuroblastoma|9500/3|Neuroblastoma
C649|Kidney|950|Neuroblastoma|9501/3|Medulloepithelioma
C649|Kidney|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C649|Kidney|950|Neuroblastoma|9503/3|Neuroepithelioma
C649|Kidney|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C649|Kidney|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C649|Kidney|959|Lymphoma|9590/3|Lymphoma
C649|Kidney|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C649|Kidney|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C649|Kidney|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C649|Kidney|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C649|Kidney|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C649|Kidney|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C649|Kidney|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C649|Kidney|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C649|Kidney|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C649|Kidney|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C649|Kidney|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C649|Kidney|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C649|Kidney|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C649|Kidney|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C649|Kidney|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C649|Kidney|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C649|Kidney|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C649|Kidney|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C649|Kidney|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C649|Kidney|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C649|Kidney|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C649|Kidney|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C649|Kidney|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C649|Kidney|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C649|Kidney|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C649|Kidney|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C649|Kidney|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C649|Kidney|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C649|Kidney|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C649|Kidney|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C649|Kidney|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C649|Kidney|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C649|Kidney|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C649|Kidney|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C649|Kidney|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C649|Kidney|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C649|Kidney|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C649|Kidney|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C649|Kidney|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C649|Kidney|973|Plasmacytoma|9731/3|Plasmacytoma
C649|Kidney|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C649|Kidney|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C649|Kidney|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C649|Kidney|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C649|Kidney|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C649|Kidney|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C649|Kidney|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C649|Kidney|975|Neoplasm|9750/3|Malignant_Histiocytosis
C649|Kidney|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C649|Kidney|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C649|Kidney|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C649|Kidney|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C649|Kidney|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C649|Kidney|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C649|Kidney|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C649|Kidney|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C649|Kidney|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C649|Kidney|981|Neoplasm|9812/3|Lymphoma
C649|Kidney|981|Neoplasm|9813/3|Lymphoma
C649|Kidney|981|Neoplasm|9814/3|Lymphoma
C649|Kidney|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C649|Kidney|981|Neoplasm|9816/3|Hypodiploid_ALL
C649|Kidney|981|Neoplasm|9817/3|Lymphoma
C649|Kidney|981|Neoplasm|9818/3|Lymphoma
C649|Kidney|981|Neoplasm|9819/3|Leukemia__B_Cell
C649|Kidney|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C649|Kidney|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C649|Kidney|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C649|Kidney|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C649|Kidney|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C649|Kidney|997|Neoplasm|9971/3|Polymorphic_PTLD
C649|Kidney|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C659, C669|Renal_Pelvis|800|Neoplasm|8000/3|Malignant_Neoplasm
C659, C669|Renal_Pelvis|800|Neoplasm|8001/3|Malignant_Cell
C659, C669|Renal_Pelvis|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C659, C669|Renal_Pelvis|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C659, C669|Renal_Pelvis|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C659, C669|Renal_Pelvis|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C659, C669|Renal_Pelvis|801|Carcinoma|8010/2|In_Situ_Cancer
C659, C669|Renal_Pelvis|801|Carcinoma|8010/3|Carcinoma
C659, C669|Renal_Pelvis|801|Carcinoma|8011/3|Malignant_Epithelioma
C659, C669|Renal_Pelvis|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C659, C669|Renal_Pelvis|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C659, C669|Renal_Pelvis|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C659, C669|Renal_Pelvis|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C659, C669|Renal_Pelvis|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C659, C669|Renal_Pelvis|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C659, C669|Renal_Pelvis|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C659, C669|Renal_Pelvis|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C659, C669|Renal_Pelvis|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C659, C669|Renal_Pelvis|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C659, C669|Renal_Pelvis|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C659, C669|Renal_Pelvis|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C659, C669|Renal_Pelvis|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C659, C669|Renal_Pelvis|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C659, C669|Renal_Pelvis|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C659, C669|Renal_Pelvis|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C659, C669|Renal_Pelvis|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C659, C669|Renal_Pelvis|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C659, C669|Renal_Pelvis|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C659, C669|Renal_Pelvis|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C659, C669|Renal_Pelvis|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C659, C669|Renal_Pelvis|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C659, C669|Renal_Pelvis|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C659, C669|Renal_Pelvis|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C659, C669|Renal_Pelvis|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C659, C669|Renal_Pelvis|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C659, C669|Renal_Pelvis|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C659, C669|Renal_Pelvis|813|Carcinoma|8130/2|Carcinoma
C659, C669|Renal_Pelvis|813|Carcinoma|8130/3|Carcinoma
C659, C669|Renal_Pelvis|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C659, C669|Renal_Pelvis|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C659, C669|Renal_Pelvis|814|Adenocarcinoma|8140/3|Adenocarcinoma
C659, C669|Renal_Pelvis|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C659, C669|Renal_Pelvis|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C659, C669|Renal_Pelvis|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C659, C669|Renal_Pelvis|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C659, C669|Renal_Pelvis|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C659, C669|Renal_Pelvis|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C659, C669|Renal_Pelvis|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C659, C669|Renal_Pelvis|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C659, C669|Renal_Pelvis|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C659, C669|Renal_Pelvis|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C659, C669|Renal_Pelvis|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C659, C669|Renal_Pelvis|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C659, C669|Renal_Pelvis|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C659, C669|Renal_Pelvis|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C659, C669|Renal_Pelvis|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C659, C669|Renal_Pelvis|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C659, C669|Renal_Pelvis|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C659, C669|Renal_Pelvis|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C659, C669|Renal_Pelvis|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C659, C669|Renal_Pelvis|880|Sarcoma|8800/3|Sarcoma
C659, C669|Renal_Pelvis|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C659, C669|Renal_Pelvis|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C659, C669|Renal_Pelvis|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C659, C669|Renal_Pelvis|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C659, C669|Renal_Pelvis|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C659, C669|Renal_Pelvis|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C659, C669|Renal_Pelvis|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C659, C669|Renal_Pelvis|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C659, C669|Renal_Pelvis|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C659, C669|Renal_Pelvis|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C659, C669|Renal_Pelvis|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C659, C669|Renal_Pelvis|882|Sarcoma|8825/3|Sarcoma
C659, C669|Renal_Pelvis|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C659, C669|Renal_Pelvis|885|Liposarcoma|8850/3|Liposarcoma
C659, C669|Renal_Pelvis|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C659, C669|Renal_Pelvis|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C659, C669|Renal_Pelvis|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C659, C669|Renal_Pelvis|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C659, C669|Renal_Pelvis|885|Liposarcoma|8855/3|Liposarcoma
C659, C669|Renal_Pelvis|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C659, C669|Renal_Pelvis|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C659, C669|Renal_Pelvis|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C659, C669|Renal_Pelvis|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C659, C669|Renal_Pelvis|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C659, C669|Renal_Pelvis|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C659, C669|Renal_Pelvis|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C659, C669|Renal_Pelvis|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C659, C669|Renal_Pelvis|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C659, C669|Renal_Pelvis|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C659, C669|Renal_Pelvis|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C659, C669|Renal_Pelvis|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C659, C669|Renal_Pelvis|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C659, C669|Renal_Pelvis|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C659, C669|Renal_Pelvis|895|Mixed_Tumor__Mullerian|8959/3|Malignant_Cystic_Nephroma
C659, C669|Renal_Pelvis|896|Nephroblastoma|8964/3|Clear_Cell_Sarcoma_Of_The_Kidney
C659, C669|Renal_Pelvis|898|Carcinosarcoma|8980/3|Carcinosarcoma
C659, C669|Renal_Pelvis|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C659, C669|Renal_Pelvis|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C659, C669|Renal_Pelvis|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C659, C669|Renal_Pelvis|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C659, C669|Renal_Pelvis|950|Neuroblastoma|9500/3|Neuroblastoma
C659, C669|Renal_Pelvis|950|Neuroblastoma|9501/3|Medulloepithelioma
C659, C669|Renal_Pelvis|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C659, C669|Renal_Pelvis|950|Neuroblastoma|9503/3|Neuroepithelioma
C659, C669|Renal_Pelvis|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C659, C669|Renal_Pelvis|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C659, C669|Renal_Pelvis|959|Lymphoma|9590/3|Lymphoma
C659, C669|Renal_Pelvis|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C659, C669|Renal_Pelvis|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C659, C669|Renal_Pelvis|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C659, C669|Renal_Pelvis|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C659, C669|Renal_Pelvis|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C659, C669|Renal_Pelvis|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C659, C669|Renal_Pelvis|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C659, C669|Renal_Pelvis|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C659, C669|Renal_Pelvis|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C659, C669|Renal_Pelvis|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C659, C669|Renal_Pelvis|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C659, C669|Renal_Pelvis|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C659, C669|Renal_Pelvis|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C659, C669|Renal_Pelvis|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C659, C669|Renal_Pelvis|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C659, C669|Renal_Pelvis|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C659, C669|Renal_Pelvis|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C659, C669|Renal_Pelvis|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C659, C669|Renal_Pelvis|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C659, C669|Renal_Pelvis|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C659, C669|Renal_Pelvis|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C659, C669|Renal_Pelvis|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C659, C669|Renal_Pelvis|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C659, C669|Renal_Pelvis|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C659, C669|Renal_Pelvis|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C659, C669|Renal_Pelvis|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C659, C669|Renal_Pelvis|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C659, C669|Renal_Pelvis|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C659, C669|Renal_Pelvis|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C659, C669|Renal_Pelvis|973|Plasmacytoma|9731/3|Plasmacytoma
C659, C669|Renal_Pelvis|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C659, C669|Renal_Pelvis|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C659, C669|Renal_Pelvis|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C659, C669|Renal_Pelvis|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C659, C669|Renal_Pelvis|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C659, C669|Renal_Pelvis|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C659, C669|Renal_Pelvis|975|Neoplasm|9750/3|Malignant_Histiocytosis
C659, C669|Renal_Pelvis|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C659, C669|Renal_Pelvis|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C659, C669|Renal_Pelvis|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C659, C669|Renal_Pelvis|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C659, C669|Renal_Pelvis|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C659, C669|Renal_Pelvis|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C659, C669|Renal_Pelvis|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C659, C669|Renal_Pelvis|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C659, C669|Renal_Pelvis|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C659, C669|Renal_Pelvis|981|Neoplasm|9812/3|Lymphoma
C659, C669|Renal_Pelvis|981|Neoplasm|9813/3|Lymphoma
C659, C669|Renal_Pelvis|981|Neoplasm|9814/3|Lymphoma
C659, C669|Renal_Pelvis|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C659, C669|Renal_Pelvis|981|Neoplasm|9816/3|Hypodiploid_ALL
C659, C669|Renal_Pelvis|981|Neoplasm|9817/3|Lymphoma
C659, C669|Renal_Pelvis|981|Neoplasm|9818/3|Lymphoma
C659, C669|Renal_Pelvis|981|Neoplasm|9819/3|Leukemia__B_Cell
C659, C669|Renal_Pelvis|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C659, C669|Renal_Pelvis|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C659, C669|Renal_Pelvis|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C659, C669|Renal_Pelvis|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C659, C669|Renal_Pelvis|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C659, C669|Renal_Pelvis|997|Neoplasm|9971/3|Polymorphic_PTLD
C659, C669|Renal_Pelvis|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C670-C679|Urinary_Bladder|800|Neoplasm|8000/3|Malignant_Neoplasm
C670-C679|Urinary_Bladder|800|Neoplasm|8001/3|Malignant_Cell
C670-C679|Urinary_Bladder|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C670-C679|Urinary_Bladder|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C670-C679|Urinary_Bladder|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C670-C679|Urinary_Bladder|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C670-C679|Urinary_Bladder|801|Carcinoma|8010/2|In_Situ_Cancer
C670-C679|Urinary_Bladder|801|Carcinoma|8010/3|Carcinoma
C670-C679|Urinary_Bladder|801|Carcinoma|8011/3|Malignant_Epithelioma
C670-C679|Urinary_Bladder|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C670-C679|Urinary_Bladder|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C670-C679|Urinary_Bladder|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C670-C679|Urinary_Bladder|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C670-C679|Urinary_Bladder|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C670-C679|Urinary_Bladder|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C670-C679|Urinary_Bladder|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C670-C679|Urinary_Bladder|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C670-C679|Urinary_Bladder|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C670-C679|Urinary_Bladder|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C670-C679|Urinary_Bladder|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C670-C679|Urinary_Bladder|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C670-C679|Urinary_Bladder|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C670-C679|Urinary_Bladder|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C670-C679|Urinary_Bladder|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C670-C679|Urinary_Bladder|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C670-C679|Urinary_Bladder|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C670-C679|Urinary_Bladder|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C670-C679|Urinary_Bladder|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C670-C679|Urinary_Bladder|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C670-C679|Urinary_Bladder|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C670-C679|Urinary_Bladder|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C670-C679|Urinary_Bladder|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C670-C679|Urinary_Bladder|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C670-C679|Urinary_Bladder|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C670-C679|Urinary_Bladder|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C670-C679|Urinary_Bladder|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C670-C679|Urinary_Bladder|813|Carcinoma|8130/2|Carcinoma
C670-C679|Urinary_Bladder|813|Carcinoma|8130/3|Carcinoma
C670-C679|Urinary_Bladder|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C670-C679|Urinary_Bladder|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C670-C679|Urinary_Bladder|814|Adenocarcinoma|8140/3|Adenocarcinoma
C670-C679|Urinary_Bladder|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C670-C679|Urinary_Bladder|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C670-C679|Urinary_Bladder|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C670-C679|Urinary_Bladder|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C670-C679|Urinary_Bladder|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C670-C679|Urinary_Bladder|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C670-C679|Urinary_Bladder|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C670-C679|Urinary_Bladder|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C670-C679|Urinary_Bladder|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C670-C679|Urinary_Bladder|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C670-C679|Urinary_Bladder|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C670-C679|Urinary_Bladder|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C670-C679|Urinary_Bladder|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C670-C679|Urinary_Bladder|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C670-C679|Urinary_Bladder|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C670-C679|Urinary_Bladder|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C670-C679|Urinary_Bladder|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C670-C679|Urinary_Bladder|857|Adenocarcinoma_With_Metaplasia|8576/3|Hepatoid_Adenocarcinoma
C670-C679|Urinary_Bladder|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C670-C679|Urinary_Bladder|880|Sarcoma|8800/3|Sarcoma
C670-C679|Urinary_Bladder|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C670-C679|Urinary_Bladder|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C670-C679|Urinary_Bladder|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C670-C679|Urinary_Bladder|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C670-C679|Urinary_Bladder|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C670-C679|Urinary_Bladder|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C670-C679|Urinary_Bladder|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C670-C679|Urinary_Bladder|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C670-C679|Urinary_Bladder|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C670-C679|Urinary_Bladder|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C670-C679|Urinary_Bladder|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C670-C679|Urinary_Bladder|882|Sarcoma|8825/3|Sarcoma
C670-C679|Urinary_Bladder|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C670-C679|Urinary_Bladder|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C670-C679|Urinary_Bladder|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C670-C679|Urinary_Bladder|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C670-C679|Urinary_Bladder|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C670-C679|Urinary_Bladder|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C670-C679|Urinary_Bladder|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C670-C679|Urinary_Bladder|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C670-C679|Urinary_Bladder|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C670-C679|Urinary_Bladder|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C670-C679|Urinary_Bladder|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C670-C679|Urinary_Bladder|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C670-C679|Urinary_Bladder|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C670-C679|Urinary_Bladder|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C670-C679|Urinary_Bladder|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C670-C679|Urinary_Bladder|898|Carcinosarcoma|8980/3|Carcinosarcoma
C670-C679|Urinary_Bladder|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C670-C679|Urinary_Bladder|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C670-C679|Urinary_Bladder|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C670-C679|Urinary_Bladder|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C670-C679|Urinary_Bladder|959|Lymphoma|9590/3|Lymphoma
C670-C679|Urinary_Bladder|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C670-C679|Urinary_Bladder|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C670-C679|Urinary_Bladder|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C670-C679|Urinary_Bladder|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C670-C679|Urinary_Bladder|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C670-C679|Urinary_Bladder|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C670-C679|Urinary_Bladder|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C670-C679|Urinary_Bladder|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C670-C679|Urinary_Bladder|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C670-C679|Urinary_Bladder|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C670-C679|Urinary_Bladder|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C670-C679|Urinary_Bladder|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C670-C679|Urinary_Bladder|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C670-C679|Urinary_Bladder|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C670-C679|Urinary_Bladder|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C670-C679|Urinary_Bladder|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C670-C679|Urinary_Bladder|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C670-C679|Urinary_Bladder|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C670-C679|Urinary_Bladder|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C670-C679|Urinary_Bladder|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C670-C679|Urinary_Bladder|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C670-C679|Urinary_Bladder|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C670-C679|Urinary_Bladder|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C670-C679|Urinary_Bladder|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C670-C679|Urinary_Bladder|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C670-C679|Urinary_Bladder|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C670-C679|Urinary_Bladder|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C670-C679|Urinary_Bladder|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C670-C679|Urinary_Bladder|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C670-C679|Urinary_Bladder|973|Plasmacytoma|9731/3|Plasmacytoma
C670-C679|Urinary_Bladder|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C670-C679|Urinary_Bladder|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C670-C679|Urinary_Bladder|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C670-C679|Urinary_Bladder|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C670-C679|Urinary_Bladder|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C670-C679|Urinary_Bladder|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C670-C679|Urinary_Bladder|975|Neoplasm|9750/3|Malignant_Histiocytosis
C670-C679|Urinary_Bladder|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C670-C679|Urinary_Bladder|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C670-C679|Urinary_Bladder|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C670-C679|Urinary_Bladder|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C670-C679|Urinary_Bladder|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C670-C679|Urinary_Bladder|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C670-C679|Urinary_Bladder|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C670-C679|Urinary_Bladder|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C670-C679|Urinary_Bladder|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C670-C679|Urinary_Bladder|981|Neoplasm|9812/3|Lymphoma
C670-C679|Urinary_Bladder|981|Neoplasm|9813/3|Lymphoma
C670-C679|Urinary_Bladder|981|Neoplasm|9814/3|Lymphoma
C670-C679|Urinary_Bladder|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C670-C679|Urinary_Bladder|981|Neoplasm|9816/3|Hypodiploid_ALL
C670-C679|Urinary_Bladder|981|Neoplasm|9817/3|Lymphoma
C670-C679|Urinary_Bladder|981|Neoplasm|9818/3|Lymphoma
C670-C679|Urinary_Bladder|981|Neoplasm|9819/3|Leukemia__B_Cell
C670-C679|Urinary_Bladder|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C670-C679|Urinary_Bladder|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C670-C679|Urinary_Bladder|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C670-C679|Urinary_Bladder|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C670-C679|Urinary_Bladder|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C670-C679|Urinary_Bladder|997|Neoplasm|9971/3|Polymorphic_PTLD
C670-C679|Urinary_Bladder|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C680-C681,C688-C689|Genitourinary_System|800|Neoplasm|8000/3|Malignant_Neoplasm
C680-C681,C688-C689|Genitourinary_System|800|Neoplasm|8001/3|Malignant_Cell
C680-C681,C688-C689|Genitourinary_System|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C680-C681,C688-C689|Genitourinary_System|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C680-C681,C688-C689|Genitourinary_System|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C680-C681,C688-C689|Genitourinary_System|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C680-C681,C688-C689|Genitourinary_System|801|Carcinoma|8010/2|In_Situ_Cancer
C680-C681,C688-C689|Genitourinary_System|801|Carcinoma|8010/3|Carcinoma
C680-C681,C688-C689|Genitourinary_System|801|Carcinoma|8011/3|Malignant_Epithelioma
C680-C681,C688-C689|Genitourinary_System|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C680-C681,C688-C689|Genitourinary_System|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C680-C681,C688-C689|Genitourinary_System|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C680-C681,C688-C689|Genitourinary_System|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C680-C681,C688-C689|Genitourinary_System|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C680-C681,C688-C689|Genitourinary_System|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C680-C681,C688-C689|Genitourinary_System|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C680-C681,C688-C689|Genitourinary_System|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C680-C681,C688-C689|Genitourinary_System|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C680-C681,C688-C689|Genitourinary_System|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C680-C681,C688-C689|Genitourinary_System|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C680-C681,C688-C689|Genitourinary_System|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C680-C681,C688-C689|Genitourinary_System|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C680-C681,C688-C689|Genitourinary_System|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C680-C681,C688-C689|Genitourinary_System|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C680-C681,C688-C689|Genitourinary_System|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C680-C681,C688-C689|Genitourinary_System|813|Carcinoma|8130/2|Carcinoma
C680-C681,C688-C689|Genitourinary_System|813|Carcinoma|8130/3|Carcinoma
C680-C681,C688-C689|Genitourinary_System|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C680-C681,C688-C689|Genitourinary_System|814|Adenocarcinoma|8140/3|Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C680-C681,C688-C689|Genitourinary_System|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C680-C681,C688-C689|Genitourinary_System|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C680-C681,C688-C689|Genitourinary_System|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C680-C681,C688-C689|Genitourinary_System|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C680-C681,C688-C689|Genitourinary_System|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C680-C681,C688-C689|Genitourinary_System|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C680-C681,C688-C689|Genitourinary_System|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C680-C681,C688-C689|Genitourinary_System|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C680-C681,C688-C689|Genitourinary_System|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C680-C681,C688-C689|Genitourinary_System|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C680-C681,C688-C689|Genitourinary_System|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C680-C681,C688-C689|Genitourinary_System|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C680-C681,C688-C689|Genitourinary_System|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C680-C681,C688-C689|Genitourinary_System|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C680-C681,C688-C689|Genitourinary_System|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C680-C681,C688-C689|Genitourinary_System|872|Melanoma|8720/3|Melanoma
C680-C681,C688-C689|Genitourinary_System|872|Melanoma|8721/3|Nodular_Melanoma
C680-C681,C688-C689|Genitourinary_System|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C680-C681,C688-C689|Genitourinary_System|872|Melanoma|8723/3|Regressing_Melanoma
C680-C681,C688-C689|Genitourinary_System|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C680-C681,C688-C689|Genitourinary_System|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C680-C681,C688-C689|Genitourinary_System|874|Nevus|8745/3|Desmoplastic_Melanoma
C680-C681,C688-C689|Genitourinary_System|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C680-C681,C688-C689|Genitourinary_System|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C680-C681,C688-C689|Genitourinary_System|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C680-C681,C688-C689|Genitourinary_System|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C680-C681,C688-C689|Genitourinary_System|880|Sarcoma|8800/3|Sarcoma
C680-C681,C688-C689|Genitourinary_System|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C680-C681,C688-C689|Genitourinary_System|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C680-C681,C688-C689|Genitourinary_System|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C680-C681,C688-C689|Genitourinary_System|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C680-C681,C688-C689|Genitourinary_System|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C680-C681,C688-C689|Genitourinary_System|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C680-C681,C688-C689|Genitourinary_System|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C680-C681,C688-C689|Genitourinary_System|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C680-C681,C688-C689|Genitourinary_System|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C680-C681,C688-C689|Genitourinary_System|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C680-C681,C688-C689|Genitourinary_System|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C680-C681,C688-C689|Genitourinary_System|882|Sarcoma|8825/3|Sarcoma
C680-C681,C688-C689|Genitourinary_System|885|Liposarcoma|8850/3|Liposarcoma
C680-C681,C688-C689|Genitourinary_System|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C680-C681,C688-C689|Genitourinary_System|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C680-C681,C688-C689|Genitourinary_System|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C680-C681,C688-C689|Genitourinary_System|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C680-C681,C688-C689|Genitourinary_System|885|Liposarcoma|8855/3|Liposarcoma
C680-C681,C688-C689|Genitourinary_System|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C680-C681,C688-C689|Genitourinary_System|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C680-C681,C688-C689|Genitourinary_System|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C680-C681,C688-C689|Genitourinary_System|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C680-C681,C688-C689|Genitourinary_System|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C680-C681,C688-C689|Genitourinary_System|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C680-C681,C688-C689|Genitourinary_System|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C680-C681,C688-C689|Genitourinary_System|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C680-C681,C688-C689|Genitourinary_System|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C680-C681,C688-C689|Genitourinary_System|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C680-C681,C688-C689|Genitourinary_System|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C680-C681,C688-C689|Genitourinary_System|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C680-C681,C688-C689|Genitourinary_System|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C680-C681,C688-C689|Genitourinary_System|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C680-C681,C688-C689|Genitourinary_System|896|Nephroblastoma|8964/3|Clear_Cell_Sarcoma_Of_The_Kidney
C680-C681,C688-C689|Genitourinary_System|898|Carcinosarcoma|8980/3|Carcinosarcoma
C680-C681,C688-C689|Genitourinary_System|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C680-C681,C688-C689|Genitourinary_System|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C680-C681,C688-C689|Genitourinary_System|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C680-C681,C688-C689|Genitourinary_System|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C680-C681,C688-C689|Genitourinary_System|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C680-C681,C688-C689|Genitourinary_System|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C680-C681,C688-C689|Genitourinary_System|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C680-C681,C688-C689|Genitourinary_System|908|Teratoma|9080/3|Immature_Teratoma
C680-C681,C688-C689|Genitourinary_System|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C680-C681,C688-C689|Genitourinary_System|908|Teratoma|9082/3|Immature_Teratoma
C680-C681,C688-C689|Genitourinary_System|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C680-C681,C688-C689|Genitourinary_System|908|Teratoma|9084/3|Teratoma
C680-C681,C688-C689|Genitourinary_System|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C680-C681,C688-C689|Genitourinary_System|911|Mesonephroma|9110/3|Mesonephroma
C680-C681,C688-C689|Genitourinary_System|950|Neuroblastoma|9500/3|Neuroblastoma
C680-C681,C688-C689|Genitourinary_System|950|Neuroblastoma|9501/3|Medulloepithelioma
C680-C681,C688-C689|Genitourinary_System|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C680-C681,C688-C689|Genitourinary_System|950|Neuroblastoma|9503/3|Neuroepithelioma
C680-C681,C688-C689|Genitourinary_System|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C680-C681,C688-C689|Genitourinary_System|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C680-C681,C688-C689|Genitourinary_System|959|Lymphoma|9590/3|Lymphoma
C680-C681,C688-C689|Genitourinary_System|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C680-C681,C688-C689|Genitourinary_System|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C680-C681,C688-C689|Genitourinary_System|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C680-C681,C688-C689|Genitourinary_System|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C680-C681,C688-C689|Genitourinary_System|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C680-C681,C688-C689|Genitourinary_System|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C680-C681,C688-C689|Genitourinary_System|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C680-C681,C688-C689|Genitourinary_System|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C680-C681,C688-C689|Genitourinary_System|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C680-C681,C688-C689|Genitourinary_System|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C680-C681,C688-C689|Genitourinary_System|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C680-C681,C688-C689|Genitourinary_System|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C680-C681,C688-C689|Genitourinary_System|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C680-C681,C688-C689|Genitourinary_System|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C680-C681,C688-C689|Genitourinary_System|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C680-C681,C688-C689|Genitourinary_System|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C680-C681,C688-C689|Genitourinary_System|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C680-C681,C688-C689|Genitourinary_System|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C680-C681,C688-C689|Genitourinary_System|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C680-C681,C688-C689|Genitourinary_System|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C680-C681,C688-C689|Genitourinary_System|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C680-C681,C688-C689|Genitourinary_System|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C680-C681,C688-C689|Genitourinary_System|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C680-C681,C688-C689|Genitourinary_System|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C680-C681,C688-C689|Genitourinary_System|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C680-C681,C688-C689|Genitourinary_System|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C680-C681,C688-C689|Genitourinary_System|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C680-C681,C688-C689|Genitourinary_System|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C680-C681,C688-C689|Genitourinary_System|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C680-C681,C688-C689|Genitourinary_System|973|Plasmacytoma|9731/3|Plasmacytoma
C680-C681,C688-C689|Genitourinary_System|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C680-C681,C688-C689|Genitourinary_System|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C680-C681,C688-C689|Genitourinary_System|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C680-C681,C688-C689|Genitourinary_System|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C680-C681,C688-C689|Genitourinary_System|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C680-C681,C688-C689|Genitourinary_System|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C680-C681,C688-C689|Genitourinary_System|975|Neoplasm|9750/3|Malignant_Histiocytosis
C680-C681,C688-C689|Genitourinary_System|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C680-C681,C688-C689|Genitourinary_System|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C680-C681,C688-C689|Genitourinary_System|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C680-C681,C688-C689|Genitourinary_System|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C680-C681,C688-C689|Genitourinary_System|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C680-C681,C688-C689|Genitourinary_System|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C680-C681,C688-C689|Genitourinary_System|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C680-C681,C688-C689|Genitourinary_System|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9812/3|Lymphoma
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9813/3|Lymphoma
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9814/3|Lymphoma
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9816/3|Hypodiploid_ALL
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9817/3|Lymphoma
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9818/3|Lymphoma
C680-C681,C688-C689|Genitourinary_System|981|Neoplasm|9819/3|Leukemia__B_Cell
C680-C681,C688-C689|Genitourinary_System|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C680-C681,C688-C689|Genitourinary_System|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C680-C681,C688-C689|Genitourinary_System|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C680-C681,C688-C689|Genitourinary_System|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C680-C681,C688-C689|Genitourinary_System|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C680-C681,C688-C689|Genitourinary_System|997|Neoplasm|9971/3|Polymorphic_PTLD
C680-C681,C688-C689|Genitourinary_System|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C690-C691, C693, C695-C698|Lacrimal_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C690-C691, C693, C695-C698|Lacrimal_Gland|800|Neoplasm|8001/3|Malignant_Cell
C690-C691, C693, C695-C698|Lacrimal_Gland|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C690-C691, C693, C695-C698|Lacrimal_Gland|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C690-C691, C693, C695-C698|Lacrimal_Gland|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C690-C691, C693, C695-C698|Lacrimal_Gland|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C690-C691, C693, C695-C698|Lacrimal_Gland|801|Carcinoma|8010/2|In_Situ_Cancer
C690-C691, C693, C695-C698|Lacrimal_Gland|801|Carcinoma|8010/3|Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|801|Carcinoma|8011/3|Malignant_Epithelioma
C690-C691, C693, C695-C698|Lacrimal_Gland|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C690-C691, C693, C695-C698|Lacrimal_Gland|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C690-C691, C693, C695-C698|Lacrimal_Gland|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|813|Carcinoma|8130/2|Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|813|Carcinoma|8130/3|Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C690-C691, C693, C695-C698|Lacrimal_Gland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C690-C691, C693, C695-C698|Lacrimal_Gland|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C690-C691, C693, C695-C698|Lacrimal_Gland|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C690-C691, C693, C695-C698|Lacrimal_Gland|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C690-C691, C693, C695-C698|Lacrimal_Gland|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|872|Melanoma|8720/3|Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|872|Melanoma|8721/3|Nodular_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|872|Melanoma|8723/3|Regressing_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C690-C691, C693, C695-C698|Lacrimal_Gland|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|874|Nevus|8745/3|Desmoplastic_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|877|Epithelioid_Cell_Melanoma|8773/3|Type_A_Spindle_Cell_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|877|Epithelioid_Cell_Melanoma|8774/3|Type_B_Spindle_Cell_Melanoma
C690-C691, C693, C695-C698|Lacrimal_Gland|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C690-C691, C693, C695-C698|Lacrimal_Gland|882|Sarcoma|8825/3|Sarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C690-C691, C693, C695-C698|Lacrimal_Gland|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C690-C691, C693, C695-C698|Lacrimal_Gland|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C690-C691, C693, C695-C698|Lacrimal_Gland|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C690-C691, C693, C695-C698|Lacrimal_Gland|959|Lymphoma|9590/3|Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C690-C691, C693, C695-C698|Lacrimal_Gland|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C690-C691, C693, C695-C698|Lacrimal_Gland|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C690-C691, C693, C695-C698|Lacrimal_Gland|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C690-C691, C693, C695-C698|Lacrimal_Gland|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C690-C691, C693, C695-C698|Lacrimal_Gland|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C690-C691, C693, C695-C698|Lacrimal_Gland|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C690-C691, C693, C695-C698|Lacrimal_Gland|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C690-C691, C693, C695-C698|Lacrimal_Gland|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C690-C691, C693, C695-C698|Lacrimal_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C690-C691, C693, C695-C698|Lacrimal_Gland|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C690-C691, C693, C695-C698|Lacrimal_Gland|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C690-C691, C693, C695-C698|Lacrimal_Gland|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C690-C691, C693, C695-C698|Lacrimal_Gland|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|973|Plasmacytoma|9731/3|Plasmacytoma
C690-C691, C693, C695-C698|Lacrimal_Gland|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C690-C691, C693, C695-C698|Lacrimal_Gland|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C690-C691, C693, C695-C698|Lacrimal_Gland|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C690-C691, C693, C695-C698|Lacrimal_Gland|975|Neoplasm|9750/3|Malignant_Histiocytosis
C690-C691, C693, C695-C698|Lacrimal_Gland|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C690-C691, C693, C695-C698|Lacrimal_Gland|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C690-C691, C693, C695-C698|Lacrimal_Gland|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C690-C691, C693, C695-C698|Lacrimal_Gland|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C690-C691, C693, C695-C698|Lacrimal_Gland|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9812/3|Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9813/3|Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9814/3|Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9816/3|Hypodiploid_ALL
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9817/3|Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9818/3|Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|981|Neoplasm|9819/3|Leukemia__B_Cell
C690-C691, C693, C695-C698|Lacrimal_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C690-C691, C693, C695-C698|Lacrimal_Gland|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C690-C691, C693, C695-C698|Lacrimal_Gland|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C690-C691, C693, C695-C698|Lacrimal_Gland|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C690-C691, C693, C695-C698|Lacrimal_Gland|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C690-C691, C693, C695-C698|Lacrimal_Gland|997|Neoplasm|9971/3|Polymorphic_PTLD
C690-C691, C693, C695-C698|Lacrimal_Gland|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C692|Retina|800|Neoplasm|8000/3|Malignant_Neoplasm
C692|Retina|800|Neoplasm|8001/3|Malignant_Cell
C692|Retina|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C692|Retina|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C692|Retina|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C692|Retina|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C692|Retina|801|Carcinoma|8010/2|In_Situ_Cancer
C692|Retina|801|Carcinoma|8010/3|Carcinoma
C692|Retina|801|Carcinoma|8011/3|Malignant_Epithelioma
C692|Retina|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C692|Retina|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C692|Retina|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C692|Retina|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C692|Retina|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C692|Retina|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C692|Retina|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C692|Retina|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C692|Retina|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C692|Retina|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C692|Retina|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C692|Retina|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C692|Retina|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C692|Retina|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C692|Retina|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C692|Retina|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C692|Retina|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C692|Retina|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C692|Retina|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C692|Retina|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C692|Retina|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C692|Retina|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C692|Retina|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C692|Retina|813|Carcinoma|8130/2|Carcinoma
C692|Retina|813|Carcinoma|8130/3|Carcinoma
C692|Retina|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C692|Retina|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C692|Retina|814|Adenocarcinoma|8140/3|Adenocarcinoma
C692|Retina|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C692|Retina|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C692|Retina|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C692|Retina|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C692|Retina|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C692|Retina|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C692|Retina|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C692|Retina|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C692|Retina|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C692|Retina|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C692|Retina|872|Melanoma|8720/3|Melanoma
C692|Retina|872|Melanoma|8721/3|Nodular_Melanoma
C692|Retina|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C692|Retina|872|Melanoma|8723/3|Regressing_Melanoma
C692|Retina|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C692|Retina|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C692|Retina|874|Nevus|8745/3|Desmoplastic_Melanoma
C692|Retina|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C692|Retina|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C692|Retina|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C692|Retina|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C692|Retina|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C692|Retina|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C692|Retina|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C692|Retina|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C692|Retina|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C692|Retina|882|Sarcoma|8825/3|Sarcoma
C692|Retina|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C692|Retina|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C692|Retina|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C692|Retina|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C692|Retina|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C692|Retina|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C692|Retina|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C692|Retina|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C692|Retina|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C692|Retina|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C692|Retina|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C692|Retina|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C692|Retina|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C692|Retina|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C692|Retina|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C692|Retina|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C692|Retina|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C692|Retina|951|Retinoblastoma|9510/3|Retinoblastoma
C692|Retina|951|Retinoblastoma|9511/3|Differentiated_Retinoblastoma
C692|Retina|951|Retinoblastoma|9512/3|Undifferentiated_Retinoblastoma
C692|Retina|951|Retinoblastoma|9513/3|Diffuse_Retinoblastoma
C692|Retina|959|Lymphoma|9590/3|Lymphoma
C692|Retina|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C692|Retina|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C692|Retina|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C692|Retina|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C692|Retina|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C692|Retina|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C692|Retina|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C692|Retina|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C692|Retina|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C692|Retina|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C692|Retina|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C692|Retina|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C692|Retina|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C692|Retina|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C692|Retina|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C692|Retina|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C692|Retina|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C692|Retina|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C692|Retina|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C692|Retina|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C692|Retina|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C692|Retina|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C692|Retina|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C692|Retina|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C692|Retina|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C692|Retina|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C692|Retina|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C692|Retina|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C692|Retina|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C692|Retina|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C692|Retina|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C692|Retina|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C692|Retina|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C692|Retina|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C692|Retina|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C692|Retina|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C692|Retina|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C692|Retina|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C692|Retina|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C692|Retina|973|Plasmacytoma|9731/3|Plasmacytoma
C692|Retina|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C692|Retina|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C692|Retina|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C692|Retina|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C692|Retina|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C692|Retina|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C692|Retina|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C692|Retina|975|Neoplasm|9750/3|Malignant_Histiocytosis
C692|Retina|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C692|Retina|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C692|Retina|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C692|Retina|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C692|Retina|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C692|Retina|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C692|Retina|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C692|Retina|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C692|Retina|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C692|Retina|981|Neoplasm|9812/3|Lymphoma
C692|Retina|981|Neoplasm|9813/3|Lymphoma
C692|Retina|981|Neoplasm|9814/3|Lymphoma
C692|Retina|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C692|Retina|981|Neoplasm|9816/3|Hypodiploid_ALL
C692|Retina|981|Neoplasm|9817/3|Lymphoma
C692|Retina|981|Neoplasm|9818/3|Lymphoma
C692|Retina|981|Neoplasm|9819/3|Leukemia__B_Cell
C692|Retina|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C692|Retina|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C692|Retina|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C692|Retina|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C692|Retina|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C692|Retina|997|Neoplasm|9971/3|Polymorphic_PTLD
C692|Retina|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C694|Eye|800|Neoplasm|8000/3|Malignant_Neoplasm
C694|Eye|800|Neoplasm|8001/3|Malignant_Cell
C694|Eye|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C694|Eye|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C694|Eye|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C694|Eye|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C694|Eye|801|Carcinoma|8010/2|In_Situ_Cancer
C694|Eye|801|Carcinoma|8010/3|Carcinoma
C694|Eye|801|Carcinoma|8011/3|Malignant_Epithelioma
C694|Eye|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C694|Eye|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C694|Eye|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C694|Eye|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C694|Eye|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C694|Eye|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C694|Eye|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C694|Eye|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C694|Eye|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C694|Eye|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C694|Eye|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C694|Eye|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C694|Eye|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C694|Eye|808|Lymphoepithelial_Carcinoma|8081/2|Bowen_Disease
C694|Eye|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C694|Eye|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C694|Eye|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C694|Eye|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C694|Eye|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C694|Eye|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C694|Eye|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C694|Eye|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C694|Eye|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C694|Eye|813|Carcinoma|8130/2|Carcinoma
C694|Eye|813|Carcinoma|8130/3|Carcinoma
C694|Eye|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C694|Eye|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C694|Eye|814|Adenocarcinoma|8140/3|Adenocarcinoma
C694|Eye|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C694|Eye|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C694|Eye|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C694|Eye|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C694|Eye|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C694|Eye|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C694|Eye|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C694|Eye|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C694|Eye|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C694|Eye|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C694|Eye|872|Melanoma|8720/3|Melanoma
C694|Eye|872|Melanoma|8721/3|Nodular_Melanoma
C694|Eye|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C694|Eye|872|Melanoma|8723/3|Regressing_Melanoma
C694|Eye|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C694|Eye|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C694|Eye|874|Nevus|8745/3|Desmoplastic_Melanoma
C694|Eye|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C694|Eye|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C694|Eye|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C694|Eye|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C694|Eye|877|Epithelioid_Cell_Melanoma|8773/3|Type_A_Spindle_Cell_Melanoma
C694|Eye|877|Epithelioid_Cell_Melanoma|8774/3|Type_B_Spindle_Cell_Melanoma
C694|Eye|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C694|Eye|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C694|Eye|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C694|Eye|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C694|Eye|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C694|Eye|882|Sarcoma|8825/3|Sarcoma
C694|Eye|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C694|Eye|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C694|Eye|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C694|Eye|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C694|Eye|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C694|Eye|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C694|Eye|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C694|Eye|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C694|Eye|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C694|Eye|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C694|Eye|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C694|Eye|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C694|Eye|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C694|Eye|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C694|Eye|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C694|Eye|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C694|Eye|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C694|Eye|959|Lymphoma|9590/3|Lymphoma
C694|Eye|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C694|Eye|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C694|Eye|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C694|Eye|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C694|Eye|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C694|Eye|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C694|Eye|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C694|Eye|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C694|Eye|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C694|Eye|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C694|Eye|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C694|Eye|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C694|Eye|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C694|Eye|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C694|Eye|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C694|Eye|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C694|Eye|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C694|Eye|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C694|Eye|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C694|Eye|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C694|Eye|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C694|Eye|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C694|Eye|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C694|Eye|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C694|Eye|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C694|Eye|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C694|Eye|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C694|Eye|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C694|Eye|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C694|Eye|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C694|Eye|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C694|Eye|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C694|Eye|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C694|Eye|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C694|Eye|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C694|Eye|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C694|Eye|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C694|Eye|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C694|Eye|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C694|Eye|973|Plasmacytoma|9731/3|Plasmacytoma
C694|Eye|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C694|Eye|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C694|Eye|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C694|Eye|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C694|Eye|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C694|Eye|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C694|Eye|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C694|Eye|975|Neoplasm|9750/3|Malignant_Histiocytosis
C694|Eye|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C694|Eye|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C694|Eye|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C694|Eye|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C694|Eye|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C694|Eye|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C694|Eye|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C694|Eye|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C694|Eye|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C694|Eye|981|Neoplasm|9812/3|Lymphoma
C694|Eye|981|Neoplasm|9813/3|Lymphoma
C694|Eye|981|Neoplasm|9814/3|Lymphoma
C694|Eye|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C694|Eye|981|Neoplasm|9816/3|Hypodiploid_ALL
C694|Eye|981|Neoplasm|9817/3|Lymphoma
C694|Eye|981|Neoplasm|9818/3|Lymphoma
C694|Eye|981|Neoplasm|9819/3|Leukemia__B_Cell
C694|Eye|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C694|Eye|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C694|Eye|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C694|Eye|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C694|Eye|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C694|Eye|997|Neoplasm|9971/3|Polymorphic_PTLD
C694|Eye|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C699|Eye|800|Neoplasm|8000/3|Malignant_Neoplasm
C699|Eye|800|Neoplasm|8001/3|Malignant_Cell
C699|Eye|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C699|Eye|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C699|Eye|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C699|Eye|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C699|Eye|801|Carcinoma|8010/2|In_Situ_Cancer
C699|Eye|801|Carcinoma|8010/3|Carcinoma
C699|Eye|801|Carcinoma|8011/3|Malignant_Epithelioma
C699|Eye|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C699|Eye|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C699|Eye|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C699|Eye|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C699|Eye|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C699|Eye|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C699|Eye|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C699|Eye|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C699|Eye|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C699|Eye|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C699|Eye|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C699|Eye|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C699|Eye|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C699|Eye|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C699|Eye|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C699|Eye|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C699|Eye|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C699|Eye|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C699|Eye|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C699|Eye|813|Carcinoma|8130/2|Carcinoma
C699|Eye|813|Carcinoma|8130/3|Carcinoma
C699|Eye|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C699|Eye|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C699|Eye|814|Adenocarcinoma|8140/3|Adenocarcinoma
C699|Eye|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C699|Eye|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C699|Eye|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C699|Eye|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C699|Eye|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C699|Eye|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C699|Eye|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C699|Eye|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C699|Eye|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C699|Eye|872|Melanoma|8720/2|Stage_0_Skin_Melanoma
C699|Eye|872|Melanoma|8720/3|Melanoma
C699|Eye|872|Melanoma|8721/3|Nodular_Melanoma
C699|Eye|872|Melanoma|8722/3|Balloon_Cell_Melanoma
C699|Eye|872|Melanoma|8723/3|Regressing_Melanoma
C699|Eye|873|Melanoma__Amelanotic|8730/3|Melanoma__Amelanotic
C699|Eye|874|Nevus|8743/3|Superficial_Spreading_Melanoma
C699|Eye|874|Nevus|8745/3|Desmoplastic_Melanoma
C699|Eye|874|Nevus|8746/3|Mucosal_Lentiginous_Melanoma
C699|Eye|877|Epithelioid_Cell_Melanoma|8770/3|Spindle_Cell_Melanoma
C699|Eye|877|Epithelioid_Cell_Melanoma|8771/3|Epithelioid_Cell_Melanoma
C699|Eye|877|Epithelioid_Cell_Melanoma|8772/3|Spindle_Cell_Melanoma
C699|Eye|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C699|Eye|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C699|Eye|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C699|Eye|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C699|Eye|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C699|Eye|882|Sarcoma|8825/3|Sarcoma
C699|Eye|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C699|Eye|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C699|Eye|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C699|Eye|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C699|Eye|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C699|Eye|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C699|Eye|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C699|Eye|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C699|Eye|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C699|Eye|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C699|Eye|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C699|Eye|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C699|Eye|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C699|Eye|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C699|Eye|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C699|Eye|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C699|Eye|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C699|Eye|951|Retinoblastoma|9510/3|Retinoblastoma
C699|Eye|951|Retinoblastoma|9511/3|Differentiated_Retinoblastoma
C699|Eye|951|Retinoblastoma|9512/3|Undifferentiated_Retinoblastoma
C699|Eye|951|Retinoblastoma|9513/3|Diffuse_Retinoblastoma
C699|Eye|959|Lymphoma|9590/3|Lymphoma
C699|Eye|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C699|Eye|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C699|Eye|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C699|Eye|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C699|Eye|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C699|Eye|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C699|Eye|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C699|Eye|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C699|Eye|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C699|Eye|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C699|Eye|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C699|Eye|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C699|Eye|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C699|Eye|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C699|Eye|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C699|Eye|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C699|Eye|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C699|Eye|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C699|Eye|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C699|Eye|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C699|Eye|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C699|Eye|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C699|Eye|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C699|Eye|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C699|Eye|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C699|Eye|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C699|Eye|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C699|Eye|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C699|Eye|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C699|Eye|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C699|Eye|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C699|Eye|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C699|Eye|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C699|Eye|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C699|Eye|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C699|Eye|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C699|Eye|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C699|Eye|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C699|Eye|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C699|Eye|973|Plasmacytoma|9731/3|Plasmacytoma
C699|Eye|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C699|Eye|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C699|Eye|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C699|Eye|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C699|Eye|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C699|Eye|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C699|Eye|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C699|Eye|975|Neoplasm|9750/3|Malignant_Histiocytosis
C699|Eye|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C699|Eye|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C699|Eye|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C699|Eye|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C699|Eye|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C699|Eye|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C699|Eye|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C699|Eye|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C699|Eye|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C699|Eye|981|Neoplasm|9812/3|Lymphoma
C699|Eye|981|Neoplasm|9813/3|Lymphoma
C699|Eye|981|Neoplasm|9814/3|Lymphoma
C699|Eye|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C699|Eye|981|Neoplasm|9816/3|Hypodiploid_ALL
C699|Eye|981|Neoplasm|9817/3|Lymphoma
C699|Eye|981|Neoplasm|9818/3|Lymphoma
C699|Eye|981|Neoplasm|9819/3|Leukemia__B_Cell
C699|Eye|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C699|Eye|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C699|Eye|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C699|Eye|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C699|Eye|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C699|Eye|997|Neoplasm|9971/3|Polymorphic_PTLD
C699|Eye|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C700-C701,C709|Meninges|800|Neoplasm|8000/0|Benign_Neoplasm
C700-C701,C709|Meninges|800|Neoplasm|8000/1|Neoplasm
C700-C701,C709|Meninges|800|Neoplasm|8000/3|Malignant_Neoplasm
C700-C701,C709|Meninges|800|Neoplasm|8001/0|Tumor_Cells__Benign
C700-C701,C709|Meninges|800|Neoplasm|8001/1|Neoplastic_Cell
C700-C701,C709|Meninges|800|Neoplasm|8001/3|Malignant_Cell
C700-C701,C709|Meninges|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C700-C701,C709|Meninges|872|Melanoma|8720/3|Melanoma
C700-C701,C709|Meninges|872|Melanoma|8728/0|Meningeal_Melanocytosis
C700-C701,C709|Meninges|872|Melanoma|8728/1|Meningeal_Melanocytoma
C700-C701,C709|Meninges|872|Melanoma|8728/3|Meningeal_Melanomatosis
C700-C701,C709|Meninges|880|Sarcoma|8800/0|Benign_Soft_Tissue_Neoplasm
C700-C701,C709|Meninges|880|Sarcoma|8800/3|Sarcoma
C700-C701,C709|Meninges|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C700-C701,C709|Meninges|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C700-C701,C709|Meninges|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C700-C701,C709|Meninges|881|Fibromatous_Neoplasm|8810/0|Fibroma
C700-C701,C709|Meninges|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C700-C701,C709|Meninges|881|Fibromatous_Neoplasm|8815/0|Solitary_Fibrous_Tumor
C700-C701,C709|Meninges|882|Sarcoma|8825/3|Sarcoma
C700-C701,C709|Meninges|885|Liposarcoma|8850/0|Lipoma
C700-C701,C709|Meninges|885|Liposarcoma|8851/0|Fibrolipoma
C700-C701,C709|Meninges|886|Angiolipoma|8861/0|Angiolipoma
C700-C701,C709|Meninges|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C700-C701,C709|Meninges|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C700-C701,C709|Meninges|908|Teratoma|9080/0|Mature_Teratoma
C700-C701,C709|Meninges|908|Teratoma|9080/1|Teratoma
C700-C701,C709|Meninges|908|Teratoma|9080/3|Immature_Teratoma
C700-C701,C709|Meninges|908|Teratoma|9084/0|Dermoid_Cyst
C700-C701,C709|Meninges|908|Teratoma|9084/3|Teratoma
C700-C701,C709|Meninges|912|Neoplasms__Vascular_Tissue|9120/0|Hemangioma
C700-C701,C709|Meninges|912|Neoplasms__Vascular_Tissue|9121/0|Hemangioma__Cavernous
C700-C701,C709|Meninges|915|Hemangiopericytoma|9150/0|Benign_Hemangiopericytoma
C700-C701,C709|Meninges|915|Hemangiopericytoma|9150/1|Hemangiopericytoma
C700-C701,C709|Meninges|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C700-C701,C709|Meninges|916|Hemangioblastoma|9161/1|Hemangioblastoma
C700-C701,C709|Meninges|924|Neoplasm|9240/3|Mesenchymal_Chondrosarcoma
C700-C701,C709|Meninges|953|Meningioma|9530/0|Meningioma
C700-C701,C709|Meninges|953|Meningioma|9530/1|Meningiomatosis
C700-C701,C709|Meninges|953|Meningioma|9530/3|Grade_III_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9531/0|Meningothelial_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9532/0|Fibrous_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9533/0|Psammomatous_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9534/0|Angiomatous_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9537/0|Transitional_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9538/1|Clear_Cell_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9538/3|Papillary_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9539/1|Atypical_Meningioma
C700-C701,C709|Meninges|953|Meningioma|9539/3|Meningeal_Sarcomatosis
C700-C701,C709|Meninges|959|Lymphoma|9590/3|Lymphoma
C700-C701,C709|Meninges|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C700-C701,C709|Meninges|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C700-C701,C709|Meninges|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C700-C701,C709|Meninges|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C700-C701,C709|Meninges|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C700-C701,C709|Meninges|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C700-C701,C709|Meninges|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C700-C701,C709|Meninges|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C700-C701,C709|Meninges|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C700-C701,C709|Meninges|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C700-C701,C709|Meninges|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C700-C701,C709|Meninges|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C700-C701,C709|Meninges|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C700-C701,C709|Meninges|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C700-C701,C709|Meninges|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C700-C701,C709|Meninges|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C700-C701,C709|Meninges|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C700-C701,C709|Meninges|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C700-C701,C709|Meninges|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C700-C701,C709|Meninges|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C700-C701,C709|Meninges|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C700-C701,C709|Meninges|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C700-C701,C709|Meninges|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C700-C701,C709|Meninges|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C700-C701,C709|Meninges|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C700-C701,C709|Meninges|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C700-C701,C709|Meninges|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C700-C701,C709|Meninges|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C700-C701,C709|Meninges|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C700-C701,C709|Meninges|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C700-C701,C709|Meninges|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C700-C701,C709|Meninges|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C700-C701,C709|Meninges|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C700-C701,C709|Meninges|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C700-C701,C709|Meninges|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C700-C701,C709|Meninges|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C700-C701,C709|Meninges|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C700-C701,C709|Meninges|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C700-C701,C709|Meninges|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C700-C701,C709|Meninges|973|Plasmacytoma|9731/3|Plasmacytoma
C700-C701,C709|Meninges|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C700-C701,C709|Meninges|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C700-C701,C709|Meninges|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C700-C701,C709|Meninges|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C700-C701,C709|Meninges|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C700-C701,C709|Meninges|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C700-C701,C709|Meninges|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C700-C701,C709|Meninges|975|Neoplasm|9750/3|Malignant_Histiocytosis
C700-C701,C709|Meninges|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C700-C701,C709|Meninges|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C700-C701,C709|Meninges|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C700-C701,C709|Meninges|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C700-C701,C709|Meninges|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C700-C701,C709|Meninges|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C700-C701,C709|Meninges|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C700-C701,C709|Meninges|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C700-C701,C709|Meninges|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C700-C701,C709|Meninges|981|Neoplasm|9812/3|Lymphoma
C700-C701,C709|Meninges|981|Neoplasm|9813/3|Lymphoma
C700-C701,C709|Meninges|981|Neoplasm|9814/3|Lymphoma
C700-C701,C709|Meninges|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C700-C701,C709|Meninges|981|Neoplasm|9816/3|Hypodiploid_ALL
C700-C701,C709|Meninges|981|Neoplasm|9817/3|Lymphoma
C700-C701,C709|Meninges|981|Neoplasm|9818/3|Lymphoma
C700-C701,C709|Meninges|981|Neoplasm|9819/3|Leukemia__B_Cell
C700-C701,C709|Meninges|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C700-C701,C709|Meninges|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C700-C701,C709|Meninges|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C700-C701,C709|Meninges|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C700-C701,C709|Meninges|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C700-C701,C709|Meninges|997|Neoplasm|9971/3|Polymorphic_PTLD
C700-C701,C709|Meninges|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8000/0|Benign_Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8000/1|Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8000/3|Malignant_Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8001/0|Tumor_Cells__Benign
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8001/1|Neoplastic_Cell
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8001/3|Malignant_Cell
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C710-C714, C717-C719, C720-C725|Cranial_Nerve|868|Paraganglioma|8680/1|Paraganglioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|872|Melanoma|8720/3|Melanoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|880|Sarcoma|8800/0|Benign_Soft_Tissue_Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|880|Sarcoma|8800/3|Sarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|881|Fibromatous_Neoplasm|8815/1|null
C710-C714, C717-C719, C720-C725|Cranial_Nerve|881|Fibromatous_Neoplasm|8815/3|Malignant_Hemangiopericytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|885|Liposarcoma|8850/0|Lipoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|885|Liposarcoma|8851/0|Fibrolipoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|906|Germ_Cell_Tumor|9064/3|Germinoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|908|Teratoma|9080/0|Mature_Teratoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|908|Teratoma|9080/1|Teratoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|908|Teratoma|9080/3|Immature_Teratoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|910|Choriocarcinoma|9100/3|Choriocarcinoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|912|Neoplasms__Vascular_Tissue|9120/0|Hemangioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|912|Neoplasms__Vascular_Tissue|9121/0|Hemangioma__Cavernous
C710-C714, C717-C719, C720-C725|Cranial_Nerve|912|Neoplasms__Vascular_Tissue|9122/0|Venous_Hemangioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|913|Hemangioendothelioma|9131/0|Capillary_Hemangioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|915|Hemangiopericytoma|9150/1|Hemangiopericytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|916|Hemangioblastoma|9161/1|Hemangioblastoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|937|Chordoma|9370/3|Chordoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|937|Chordoma|9371/3|Chondroid_Chordoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|938|Glioma|9380/3|Malignant_Glioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|938|Glioma|9381/3|Gliomatosis_Cerebri
C710-C714, C717-C719, C720-C725|Cranial_Nerve|938|Glioma|9382/3|Mixed_Glioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|938|Glioma|9383/1|Subependymal_Glioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|938|Glioma|9384/1|Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|938|Glioma|9385/3|Glioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|939|Ependymoma|9391/3|Ependymoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|939|Ependymoma|9392/3|Anaplastic_Ependymoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|939|Ependymoma|9393/3|Papillary_Ependymoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|939|Ependymoma|9394/1|Myxopapillary_Ependymoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|939|Ependymoma|9396/3|Ependymoma__RELA_Fusion_Positive
C710-C714, C717-C719, C720-C725|Cranial_Nerve|940|Astrocytoma|9400/3|Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|940|Astrocytoma|9401/3|Anaplastic_Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|941|Protoplasmic_Astrocytoma|9410/3|Protoplasmic_Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|941|Protoplasmic_Astrocytoma|9411/3|Gemistocytic_Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|941|Protoplasmic_Astrocytoma|9412/1|Desmoplastic_Infantile_Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|941|Protoplasmic_Astrocytoma|9413/0|Dysembryoplastic_Neuroepithelial_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|942|Fibrillary_Astrocytoma|9420/3|Fibrillary_Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|942|Fibrillary_Astrocytoma|9421/1|Pilocytic_Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|942|Fibrillary_Astrocytoma|9421/3|Pilocytic_Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|942|Fibrillary_Astrocytoma|9423/3|Polar_Spongioblastoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|942|Fibrillary_Astrocytoma|9424/3|Pleomorphic_Xanthoastrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|942|Fibrillary_Astrocytoma|9425/3|Pilomyxoid_Astrocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|943|Astroblastoma|9430/3|Astroblastoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|943|Astroblastoma|9431/1|Angiocentric_Glioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|944|Glioblastoma|9440/3|Glioblastoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|944|Glioblastoma|9441/3|Giant_Cell_Glioblastoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|944|Glioblastoma|9442/1|Gliofibroma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|944|Glioblastoma|9442/3|Gliosarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|944|Glioblastoma|9444/1|Chordoid_Glioma_Of_The_Third_Ventricle
C710-C714, C717-C719, C720-C725|Cranial_Nerve|944|Glioblastoma|9445/3|Glioblastoma__IDH_Mutant
C710-C714, C717-C719, C720-C725|Cranial_Nerve|945|Adult_Oligodendroglioma|9450/3|Adult_Oligodendroglioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|945|Adult_Oligodendroglioma|9451/3|Anaplastic_Oligodendroglioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|946|Oligodendroblastoma|9460/3|Oligodendroblastoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|947|Medulloblastoma|9473/3|Primitive_Neuroectodermal_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|947|Medulloblastoma|9475/3|Medulloblastoma__WNT_Activated
C710-C714, C717-C719, C720-C725|Cranial_Nerve|947|Medulloblastoma|9476/3|Medulloblastoma__SHH_Activated
C710-C714, C717-C719, C720-C725|Cranial_Nerve|947|Medulloblastoma|9477/3|Medulloblastoma__Non_WNT_Non_SHH
C710-C714, C717-C719, C720-C725|Cranial_Nerve|947|Medulloblastoma|9478/3|Embryonal_Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|949|Ganglioneuroblastoma|9490/0|Ganglioneuroma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|949|Ganglioneuroblastoma|9492/0|Gangliocytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9500/3|Neuroblastoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9501/3|Medulloepithelioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9503/3|Neuroepithelioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9505/0|Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9505/1|Ganglioglioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9508/3|Atypical_Teratoid_Rhabdoid_Tumor_CL372028
C710-C714, C717-C719, C720-C725|Cranial_Nerve|950|Neuroblastoma|9509/1|Papillary_Glioneuronal_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/0|Neurofibroma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/1|Neurofibromatosis
C710-C714, C717-C719, C720-C725|Cranial_Nerve|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9541/0|Melanotic_Neurofibroma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|955|Plexiform_Neurofibroma|9550/0|Plexiform_Neurofibroma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|956|Schwannoma|9560/0|Schwannoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|956|Schwannoma|9560/1|Melanotic_Schwannoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|956|Schwannoma|9562/0|Neurothekeoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|957|Perineurioma|9570/0|Neuroma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|957|Perineurioma|9571/0|Perineurioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|957|Perineurioma|9571/3|Malignant_Perineurioma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|959|Lymphoma|9590/3|Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C710-C714, C717-C719, C720-C725|Cranial_Nerve|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C710-C714, C717-C719, C720-C725|Cranial_Nerve|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C710-C714, C717-C719, C720-C725|Cranial_Nerve|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C710-C714, C717-C719, C720-C725|Cranial_Nerve|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C710-C714, C717-C719, C720-C725|Cranial_Nerve|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C710-C714, C717-C719, C720-C725|Cranial_Nerve|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C710-C714, C717-C719, C720-C725|Cranial_Nerve|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|973|Plasmacytoma|9731/3|Plasmacytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C710-C714, C717-C719, C720-C725|Cranial_Nerve|975|Neoplasm|9750/3|Malignant_Histiocytosis
C710-C714, C717-C719, C720-C725|Cranial_Nerve|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C710-C714, C717-C719, C720-C725|Cranial_Nerve|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C710-C714, C717-C719, C720-C725|Cranial_Nerve|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C710-C714, C717-C719, C720-C725|Cranial_Nerve|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9812/3|Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9813/3|Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9814/3|Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9816/3|Hypodiploid_ALL
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9817/3|Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9818/3|Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|981|Neoplasm|9819/3|Leukemia__B_Cell
C710-C714, C717-C719, C720-C725|Cranial_Nerve|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C710-C714, C717-C719, C720-C725|Cranial_Nerve|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C710-C714, C717-C719, C720-C725|Cranial_Nerve|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|993|Myeloid_Sarcoma|9930/3|Myeloid_Sarcoma
C710-C714, C717-C719, C720-C725|Cranial_Nerve|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C710-C714, C717-C719, C720-C725|Cranial_Nerve|997|Neoplasm|9971/3|Polymorphic_PTLD
C710-C714, C717-C719, C720-C725|Cranial_Nerve|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C715|Heart_Ventricle|800|Neoplasm|8000/0|Benign_Neoplasm
C715|Heart_Ventricle|800|Neoplasm|8000/1|Neoplasm
C715|Heart_Ventricle|800|Neoplasm|8000/3|Malignant_Neoplasm
C715|Heart_Ventricle|800|Neoplasm|8001/0|Tumor_Cells__Benign
C715|Heart_Ventricle|800|Neoplasm|8001/1|Neoplastic_Cell
C715|Heart_Ventricle|800|Neoplasm|8001/3|Malignant_Cell
C715|Heart_Ventricle|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C715|Heart_Ventricle|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C715|Heart_Ventricle|937|Chordoma|9370/3|Chordoma
C715|Heart_Ventricle|937|Chordoma|9371/3|Chondroid_Chordoma
C715|Heart_Ventricle|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C715|Heart_Ventricle|938|Glioma|9380/3|Malignant_Glioma
C715|Heart_Ventricle|938|Glioma|9381/3|Gliomatosis_Cerebri
C715|Heart_Ventricle|938|Glioma|9382/3|Mixed_Glioma
C715|Heart_Ventricle|938|Glioma|9383/1|Subependymal_Glioma
C715|Heart_Ventricle|938|Glioma|9384/1|Astrocytoma
C715|Heart_Ventricle|938|Glioma|9385/3|Glioma
C715|Heart_Ventricle|939|Ependymoma|9390/0|Choroid_Plexus_Papilloma
C715|Heart_Ventricle|939|Ependymoma|9390/1|Atypical_Choroid_Plexus_Papilloma
C715|Heart_Ventricle|939|Ependymoma|9390/3|Choroid_Plexus_Carcinoma
C715|Heart_Ventricle|939|Ependymoma|9391/3|Ependymoma
C715|Heart_Ventricle|939|Ependymoma|9392/3|Anaplastic_Ependymoma
C715|Heart_Ventricle|939|Ependymoma|9393/3|Papillary_Ependymoma
C715|Heart_Ventricle|939|Ependymoma|9396/3|Ependymoma__RELA_Fusion_Positive
C715|Heart_Ventricle|940|Astrocytoma|9400/3|Astrocytoma
C715|Heart_Ventricle|940|Astrocytoma|9401/3|Anaplastic_Astrocytoma
C715|Heart_Ventricle|941|Protoplasmic_Astrocytoma|9410/3|Protoplasmic_Astrocytoma
C715|Heart_Ventricle|941|Protoplasmic_Astrocytoma|9411/3|Gemistocytic_Astrocytoma
C715|Heart_Ventricle|942|Fibrillary_Astrocytoma|9420/3|Fibrillary_Astrocytoma
C715|Heart_Ventricle|942|Fibrillary_Astrocytoma|9421/1|Pilocytic_Astrocytoma
C715|Heart_Ventricle|942|Fibrillary_Astrocytoma|9421/3|Pilocytic_Astrocytoma
C715|Heart_Ventricle|942|Fibrillary_Astrocytoma|9423/3|Polar_Spongioblastoma
C715|Heart_Ventricle|942|Fibrillary_Astrocytoma|9424/3|Pleomorphic_Xanthoastrocytoma
C715|Heart_Ventricle|942|Fibrillary_Astrocytoma|9425/3|Pilomyxoid_Astrocytoma
C715|Heart_Ventricle|943|Astroblastoma|9430/3|Astroblastoma
C715|Heart_Ventricle|943|Astroblastoma|9431/1|Angiocentric_Glioma
C715|Heart_Ventricle|944|Glioblastoma|9440/3|Glioblastoma
C715|Heart_Ventricle|944|Glioblastoma|9441/3|Giant_Cell_Glioblastoma
C715|Heart_Ventricle|944|Glioblastoma|9442/3|Gliosarcoma
C715|Heart_Ventricle|944|Glioblastoma|9444/1|Chordoid_Glioma_Of_The_Third_Ventricle
C715|Heart_Ventricle|944|Glioblastoma|9445/3|Glioblastoma__IDH_Mutant
C715|Heart_Ventricle|945|Adult_Oligodendroglioma|9450/3|Adult_Oligodendroglioma
C715|Heart_Ventricle|945|Adult_Oligodendroglioma|9451/3|Anaplastic_Oligodendroglioma
C715|Heart_Ventricle|947|Medulloblastoma|9473/3|Primitive_Neuroectodermal_Tumor
C715|Heart_Ventricle|947|Medulloblastoma|9475/3|Medulloblastoma__WNT_Activated
C715|Heart_Ventricle|947|Medulloblastoma|9476/3|Medulloblastoma__SHH_Activated
C715|Heart_Ventricle|947|Medulloblastoma|9477/3|Medulloblastoma__Non_WNT_Non_SHH
C715|Heart_Ventricle|947|Medulloblastoma|9478/3|Embryonal_Neoplasm
C715|Heart_Ventricle|949|Ganglioneuroblastoma|9490/0|Ganglioneuroma
C715|Heart_Ventricle|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C715|Heart_Ventricle|949|Ganglioneuroblastoma|9492/0|Gangliocytoma
C715|Heart_Ventricle|950|Neuroblastoma|9500/3|Neuroblastoma
C715|Heart_Ventricle|950|Neuroblastoma|9501/3|Medulloepithelioma
C715|Heart_Ventricle|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C715|Heart_Ventricle|950|Neuroblastoma|9503/3|Neuroepithelioma
C715|Heart_Ventricle|950|Neuroblastoma|9505/1|Ganglioglioma
C715|Heart_Ventricle|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C715|Heart_Ventricle|950|Neuroblastoma|9506/1|Neurocytoma
C715|Heart_Ventricle|950|Neuroblastoma|9508/3|Atypical_Teratoid_Rhabdoid_Tumor_CL372028
C715|Heart_Ventricle|950|Neuroblastoma|9509/1|Papillary_Glioneuronal_Tumor
C715|Heart_Ventricle|959|Lymphoma|9590/3|Lymphoma
C715|Heart_Ventricle|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C715|Heart_Ventricle|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C715|Heart_Ventricle|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C715|Heart_Ventricle|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C715|Heart_Ventricle|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C715|Heart_Ventricle|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C715|Heart_Ventricle|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C715|Heart_Ventricle|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C715|Heart_Ventricle|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C715|Heart_Ventricle|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C715|Heart_Ventricle|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C715|Heart_Ventricle|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C715|Heart_Ventricle|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C715|Heart_Ventricle|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C715|Heart_Ventricle|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C715|Heart_Ventricle|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C715|Heart_Ventricle|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C715|Heart_Ventricle|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C715|Heart_Ventricle|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C715|Heart_Ventricle|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C715|Heart_Ventricle|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C715|Heart_Ventricle|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C715|Heart_Ventricle|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C715|Heart_Ventricle|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C715|Heart_Ventricle|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C715|Heart_Ventricle|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C715|Heart_Ventricle|973|Plasmacytoma|9731/3|Plasmacytoma
C715|Heart_Ventricle|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C715|Heart_Ventricle|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C715|Heart_Ventricle|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C715|Heart_Ventricle|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C715|Heart_Ventricle|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C715|Heart_Ventricle|975|Neoplasm|9750/3|Malignant_Histiocytosis
C715|Heart_Ventricle|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C715|Heart_Ventricle|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C715|Heart_Ventricle|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C715|Heart_Ventricle|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C715|Heart_Ventricle|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C715|Heart_Ventricle|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C715|Heart_Ventricle|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C715|Heart_Ventricle|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C715|Heart_Ventricle|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C715|Heart_Ventricle|981|Neoplasm|9812/3|Lymphoma
C715|Heart_Ventricle|981|Neoplasm|9813/3|Lymphoma
C715|Heart_Ventricle|981|Neoplasm|9814/3|Lymphoma
C715|Heart_Ventricle|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C715|Heart_Ventricle|981|Neoplasm|9816/3|Hypodiploid_ALL
C715|Heart_Ventricle|981|Neoplasm|9817/3|Lymphoma
C715|Heart_Ventricle|981|Neoplasm|9818/3|Lymphoma
C715|Heart_Ventricle|981|Neoplasm|9819/3|Leukemia__B_Cell
C715|Heart_Ventricle|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C715|Heart_Ventricle|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C715|Heart_Ventricle|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C715|Heart_Ventricle|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C715|Heart_Ventricle|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C715|Heart_Ventricle|997|Neoplasm|9971/3|Polymorphic_PTLD
C715|Heart_Ventricle|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C716|Cerebellum|800|Neoplasm|8000/0|Benign_Neoplasm
C716|Cerebellum|800|Neoplasm|8000/1|Neoplasm
C716|Cerebellum|800|Neoplasm|8000/3|Malignant_Neoplasm
C716|Cerebellum|800|Neoplasm|8001/0|Tumor_Cells__Benign
C716|Cerebellum|800|Neoplasm|8001/1|Neoplastic_Cell
C716|Cerebellum|800|Neoplasm|8001/3|Malignant_Cell
C716|Cerebellum|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C716|Cerebellum|880|Sarcoma|8800/0|Benign_Soft_Tissue_Neoplasm
C716|Cerebellum|880|Sarcoma|8800/3|Sarcoma
C716|Cerebellum|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C716|Cerebellum|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C716|Cerebellum|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C716|Cerebellum|881|Fibromatous_Neoplasm|8815/0|Solitary_Fibrous_Tumor
C716|Cerebellum|882|Sarcoma|8825/3|Sarcoma
C716|Cerebellum|885|Liposarcoma|8850/0|Lipoma
C716|Cerebellum|908|Teratoma|9080/0|Mature_Teratoma
C716|Cerebellum|908|Teratoma|9080/1|Teratoma
C716|Cerebellum|908|Teratoma|9080/3|Immature_Teratoma
C716|Cerebellum|908|Teratoma|9084/0|Dermoid_Cyst
C716|Cerebellum|912|Neoplasms__Vascular_Tissue|9120/0|Hemangioma
C716|Cerebellum|913|Hemangioendothelioma|9131/0|Capillary_Hemangioma
C716|Cerebellum|915|Hemangiopericytoma|9150/1|Hemangiopericytoma
C716|Cerebellum|916|Hemangioblastoma|9161/1|Hemangioblastoma
C716|Cerebellum|937|Chordoma|9370/3|Chordoma
C716|Cerebellum|937|Chordoma|9371/3|Chondroid_Chordoma
C716|Cerebellum|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C716|Cerebellum|938|Glioma|9380/3|Malignant_Glioma
C716|Cerebellum|938|Glioma|9381/3|Gliomatosis_Cerebri
C716|Cerebellum|938|Glioma|9382/3|Mixed_Glioma
C716|Cerebellum|938|Glioma|9383/1|Subependymal_Glioma
C716|Cerebellum|938|Glioma|9385/3|Glioma
C716|Cerebellum|939|Ependymoma|9391/3|Ependymoma
C716|Cerebellum|939|Ependymoma|9392/3|Anaplastic_Ependymoma
C716|Cerebellum|939|Ependymoma|9393/3|Papillary_Ependymoma
C716|Cerebellum|939|Ependymoma|9396/3|Ependymoma__RELA_Fusion_Positive
C716|Cerebellum|940|Astrocytoma|9400/3|Astrocytoma
C716|Cerebellum|940|Astrocytoma|9401/3|Anaplastic_Astrocytoma
C716|Cerebellum|941|Protoplasmic_Astrocytoma|9410/3|Protoplasmic_Astrocytoma
C716|Cerebellum|941|Protoplasmic_Astrocytoma|9411/3|Gemistocytic_Astrocytoma
C716|Cerebellum|942|Fibrillary_Astrocytoma|9420/3|Fibrillary_Astrocytoma
C716|Cerebellum|942|Fibrillary_Astrocytoma|9421/1|Pilocytic_Astrocytoma
C716|Cerebellum|942|Fibrillary_Astrocytoma|9421/3|Pilocytic_Astrocytoma
C716|Cerebellum|942|Fibrillary_Astrocytoma|9424/3|Pleomorphic_Xanthoastrocytoma
C716|Cerebellum|942|Fibrillary_Astrocytoma|9425/3|Pilomyxoid_Astrocytoma
C716|Cerebellum|943|Astroblastoma|9430/3|Astroblastoma
C716|Cerebellum|943|Astroblastoma|9431/1|Angiocentric_Glioma
C716|Cerebellum|944|Glioblastoma|9440/3|Glioblastoma
C716|Cerebellum|944|Glioblastoma|9441/3|Giant_Cell_Glioblastoma
C716|Cerebellum|944|Glioblastoma|9442/3|Gliosarcoma
C716|Cerebellum|944|Glioblastoma|9445/3|Glioblastoma__IDH_Mutant
C716|Cerebellum|945|Adult_Oligodendroglioma|9450/3|Adult_Oligodendroglioma
C716|Cerebellum|945|Adult_Oligodendroglioma|9451/3|Anaplastic_Oligodendroglioma
C716|Cerebellum|947|Medulloblastoma|9470/3|Medulloblastoma
C716|Cerebellum|947|Medulloblastoma|9471/3|Desmoplastic_Nodular_Medulloblastoma
C716|Cerebellum|947|Medulloblastoma|9472/3|Medullomyoblastoma
C716|Cerebellum|947|Medulloblastoma|9473/3|Primitive_Neuroectodermal_Tumor
C716|Cerebellum|947|Medulloblastoma|9474/3|Large_Cell_Medulloblastoma
C716|Cerebellum|947|Medulloblastoma|9475/3|Medulloblastoma__WNT_Activated
C716|Cerebellum|947|Medulloblastoma|9476/3|Medulloblastoma__SHH_Activated
C716|Cerebellum|947|Medulloblastoma|9477/3|Medulloblastoma__Non_WNT_Non_SHH
C716|Cerebellum|947|Medulloblastoma|9478/3|Embryonal_Neoplasm
C716|Cerebellum|948|Cerebellar_Sarcoma|9480/3|Cerebellar_Sarcoma
C716|Cerebellum|949|Ganglioneuroblastoma|9490/0|Ganglioneuroma
C716|Cerebellum|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C716|Cerebellum|949|Ganglioneuroblastoma|9492/0|Gangliocytoma
C716|Cerebellum|949|Ganglioneuroblastoma|9493/0|Lhermitte_Duclos_Disease
C716|Cerebellum|950|Neuroblastoma|9500/3|Neuroblastoma
C716|Cerebellum|950|Neuroblastoma|9501/3|Medulloepithelioma
C716|Cerebellum|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C716|Cerebellum|950|Neuroblastoma|9503/3|Neuroepithelioma
C716|Cerebellum|950|Neuroblastoma|9505/1|Ganglioglioma
C716|Cerebellum|950|Neuroblastoma|9506/1|Neurocytoma
C716|Cerebellum|950|Neuroblastoma|9508/3|Atypical_Teratoid_Rhabdoid_Tumor_CL372028
C716|Cerebellum|950|Neuroblastoma|9509/1|Papillary_Glioneuronal_Tumor
C716|Cerebellum|959|Lymphoma|9590/3|Lymphoma
C716|Cerebellum|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C716|Cerebellum|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C716|Cerebellum|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C716|Cerebellum|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C716|Cerebellum|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C716|Cerebellum|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C716|Cerebellum|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C716|Cerebellum|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C716|Cerebellum|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C716|Cerebellum|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C716|Cerebellum|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C716|Cerebellum|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C716|Cerebellum|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C716|Cerebellum|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C716|Cerebellum|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C716|Cerebellum|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C716|Cerebellum|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C716|Cerebellum|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C716|Cerebellum|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C716|Cerebellum|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C716|Cerebellum|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C716|Cerebellum|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C716|Cerebellum|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C716|Cerebellum|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C716|Cerebellum|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C716|Cerebellum|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C716|Cerebellum|973|Plasmacytoma|9731/3|Plasmacytoma
C716|Cerebellum|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C716|Cerebellum|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C716|Cerebellum|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C716|Cerebellum|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C716|Cerebellum|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C716|Cerebellum|975|Neoplasm|9750/3|Malignant_Histiocytosis
C716|Cerebellum|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C716|Cerebellum|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C716|Cerebellum|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C716|Cerebellum|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C716|Cerebellum|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C716|Cerebellum|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C716|Cerebellum|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C716|Cerebellum|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C716|Cerebellum|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C716|Cerebellum|981|Neoplasm|9812/3|Lymphoma
C716|Cerebellum|981|Neoplasm|9813/3|Lymphoma
C716|Cerebellum|981|Neoplasm|9814/3|Lymphoma
C716|Cerebellum|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C716|Cerebellum|981|Neoplasm|9816/3|Hypodiploid_ALL
C716|Cerebellum|981|Neoplasm|9817/3|Lymphoma
C716|Cerebellum|981|Neoplasm|9818/3|Lymphoma
C716|Cerebellum|981|Neoplasm|9819/3|Leukemia__B_Cell
C716|Cerebellum|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C716|Cerebellum|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C716|Cerebellum|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C716|Cerebellum|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C716|Cerebellum|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C716|Cerebellum|997|Neoplasm|9971/3|Polymorphic_PTLD
C716|Cerebellum|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C728-C729|Central_Nervous_System|800|Neoplasm|8000/0|Benign_Neoplasm
C728-C729|Central_Nervous_System|800|Neoplasm|8000/1|Neoplasm
C728-C729|Central_Nervous_System|800|Neoplasm|8000/3|Malignant_Neoplasm
C728-C729|Central_Nervous_System|800|Neoplasm|8001/0|Tumor_Cells__Benign
C728-C729|Central_Nervous_System|800|Neoplasm|8001/1|Neoplastic_Cell
C728-C729|Central_Nervous_System|800|Neoplasm|8001/3|Malignant_Cell
C728-C729|Central_Nervous_System|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C728-C729|Central_Nervous_System|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C728-C729|Central_Nervous_System|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C728-C729|Central_Nervous_System|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C728-C729|Central_Nervous_System|880|Sarcoma|8800/0|Benign_Soft_Tissue_Neoplasm
C728-C729|Central_Nervous_System|880|Sarcoma|8800/3|Sarcoma
C728-C729|Central_Nervous_System|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C728-C729|Central_Nervous_System|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C728-C729|Central_Nervous_System|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C728-C729|Central_Nervous_System|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C728-C729|Central_Nervous_System|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C728-C729|Central_Nervous_System|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C728-C729|Central_Nervous_System|885|Liposarcoma|8850/0|Lipoma
C728-C729|Central_Nervous_System|885|Liposarcoma|8850/1|Atypical_Lipoma
C728-C729|Central_Nervous_System|885|Liposarcoma|8850/3|Liposarcoma
C728-C729|Central_Nervous_System|886|Angiolipoma|8861/0|Angiolipoma
C728-C729|Central_Nervous_System|889|Myomatous_Neoplasm|8890/0|Fibroid_Tumor
C728-C729|Central_Nervous_System|889|Myomatous_Neoplasm|8890/1|Leiomyomatosis
C728-C729|Central_Nervous_System|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C728-C729|Central_Nervous_System|889|Myomatous_Neoplasm|8897/1|Smooth_Muscle_Neoplasm
C728-C729|Central_Nervous_System|890|Rhabdomyosarcoma|8900/0|Rhabdomyoma
C728-C729|Central_Nervous_System|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C728-C729|Central_Nervous_System|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C728-C729|Central_Nervous_System|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C728-C729|Central_Nervous_System|906|Germ_Cell_Tumor|9064/3|Germinoma
C728-C729|Central_Nervous_System|908|Teratoma|9080/1|Teratoma
C728-C729|Central_Nervous_System|908|Teratoma|9080/3|Immature_Teratoma
C728-C729|Central_Nervous_System|908|Teratoma|9082/3|Immature_Teratoma
C728-C729|Central_Nervous_System|908|Teratoma|9084/0|Dermoid_Cyst
C728-C729|Central_Nervous_System|908|Teratoma|9084/3|Teratoma
C728-C729|Central_Nervous_System|912|Neoplasms__Vascular_Tissue|9120/0|Hemangioma
C728-C729|Central_Nervous_System|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C728-C729|Central_Nervous_System|912|Neoplasms__Vascular_Tissue|9121/0|Hemangioma__Cavernous
C728-C729|Central_Nervous_System|913|Hemangioendothelioma|9130/0|Benign_Hemangioendothelioma
C728-C729|Central_Nervous_System|913|Hemangioendothelioma|9130/1|Hemangioendothelioma
C728-C729|Central_Nervous_System|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C728-C729|Central_Nervous_System|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C728-C729|Central_Nervous_System|915|Hemangiopericytoma|9150/0|Benign_Hemangiopericytoma
C728-C729|Central_Nervous_System|915|Hemangiopericytoma|9150/1|Hemangiopericytoma
C728-C729|Central_Nervous_System|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C728-C729|Central_Nervous_System|916|Hemangioblastoma|9161/1|Hemangioblastoma
C728-C729|Central_Nervous_System|926|Ewing_Sarcoma|9260/3|Ewing_Sarcoma
C728-C729|Central_Nervous_System|937|Chordoma|9370/3|Chordoma
C728-C729|Central_Nervous_System|937|Chordoma|9371/3|Chondroid_Chordoma
C728-C729|Central_Nervous_System|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C728-C729|Central_Nervous_System|950|Neuroblastoma|9500/3|Neuroblastoma
C728-C729|Central_Nervous_System|950|Neuroblastoma|9501/3|Medulloepithelioma
C728-C729|Central_Nervous_System|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C728-C729|Central_Nervous_System|950|Neuroblastoma|9503/3|Neuroepithelioma
C728-C729|Central_Nervous_System|950|Neuroblastoma|9508/3|Atypical_Teratoid_Rhabdoid_Tumor_CL372028
C728-C729|Central_Nervous_System|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/0|Neurofibroma
C728-C729|Central_Nervous_System|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/1|Neurofibromatosis
C728-C729|Central_Nervous_System|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C728-C729|Central_Nervous_System|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9541/0|Melanotic_Neurofibroma
C728-C729|Central_Nervous_System|955|Plexiform_Neurofibroma|9550/0|Plexiform_Neurofibroma
C728-C729|Central_Nervous_System|956|Schwannoma|9560/0|Schwannoma
C728-C729|Central_Nervous_System|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C728-C729|Central_Nervous_System|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C728-C729|Central_Nervous_System|956|Schwannoma|9562/0|Neurothekeoma
C728-C729|Central_Nervous_System|957|Perineurioma|9570/0|Neuroma
C728-C729|Central_Nervous_System|957|Perineurioma|9571/0|Perineurioma
C728-C729|Central_Nervous_System|957|Perineurioma|9571/3|Malignant_Perineurioma
C728-C729|Central_Nervous_System|959|Lymphoma|9590/3|Lymphoma
C728-C729|Central_Nervous_System|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C728-C729|Central_Nervous_System|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C728-C729|Central_Nervous_System|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C728-C729|Central_Nervous_System|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C728-C729|Central_Nervous_System|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C728-C729|Central_Nervous_System|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C728-C729|Central_Nervous_System|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C728-C729|Central_Nervous_System|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C728-C729|Central_Nervous_System|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C728-C729|Central_Nervous_System|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C728-C729|Central_Nervous_System|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C728-C729|Central_Nervous_System|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C728-C729|Central_Nervous_System|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C728-C729|Central_Nervous_System|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C728-C729|Central_Nervous_System|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C728-C729|Central_Nervous_System|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C728-C729|Central_Nervous_System|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C728-C729|Central_Nervous_System|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C728-C729|Central_Nervous_System|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C728-C729|Central_Nervous_System|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C728-C729|Central_Nervous_System|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C728-C729|Central_Nervous_System|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C728-C729|Central_Nervous_System|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C728-C729|Central_Nervous_System|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C728-C729|Central_Nervous_System|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C728-C729|Central_Nervous_System|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C728-C729|Central_Nervous_System|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C728-C729|Central_Nervous_System|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C728-C729|Central_Nervous_System|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C728-C729|Central_Nervous_System|973|Plasmacytoma|9731/3|Plasmacytoma
C728-C729|Central_Nervous_System|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C728-C729|Central_Nervous_System|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C728-C729|Central_Nervous_System|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C728-C729|Central_Nervous_System|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C728-C729|Central_Nervous_System|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C728-C729|Central_Nervous_System|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C728-C729|Central_Nervous_System|975|Neoplasm|9750/3|Malignant_Histiocytosis
C728-C729|Central_Nervous_System|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C728-C729|Central_Nervous_System|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C728-C729|Central_Nervous_System|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C728-C729|Central_Nervous_System|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C728-C729|Central_Nervous_System|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C728-C729|Central_Nervous_System|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C728-C729|Central_Nervous_System|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C728-C729|Central_Nervous_System|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C728-C729|Central_Nervous_System|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C728-C729|Central_Nervous_System|981|Neoplasm|9812/3|Lymphoma
C728-C729|Central_Nervous_System|981|Neoplasm|9813/3|Lymphoma
C728-C729|Central_Nervous_System|981|Neoplasm|9814/3|Lymphoma
C728-C729|Central_Nervous_System|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C728-C729|Central_Nervous_System|981|Neoplasm|9816/3|Hypodiploid_ALL
C728-C729|Central_Nervous_System|981|Neoplasm|9817/3|Lymphoma
C728-C729|Central_Nervous_System|981|Neoplasm|9818/3|Lymphoma
C728-C729|Central_Nervous_System|981|Neoplasm|9819/3|Leukemia__B_Cell
C728-C729|Central_Nervous_System|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C728-C729|Central_Nervous_System|982|Lymphoid_Leukemia|9827/3|Adult_T_cell_Leukemia
C728-C729|Central_Nervous_System|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C728-C729|Central_Nervous_System|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C728-C729|Central_Nervous_System|986|Myeloid_Leukemia|9861/3|Acute_Myeloid_Leukemia
C728-C729|Central_Nervous_System|993|Myeloid_Sarcoma|9930/3|Myeloid_Sarcoma
C728-C729|Central_Nervous_System|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C728-C729|Central_Nervous_System|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C728-C729|Central_Nervous_System|997|Neoplasm|9971/3|Polymorphic_PTLD
C728-C729|Central_Nervous_System|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C739|Thyroid_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C739|Thyroid_Gland|800|Neoplasm|8001/3|Malignant_Cell
C739|Thyroid_Gland|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C739|Thyroid_Gland|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C739|Thyroid_Gland|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C739|Thyroid_Gland|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C739|Thyroid_Gland|801|Carcinoma|8010/2|In_Situ_Cancer
C739|Thyroid_Gland|801|Carcinoma|8010/3|Carcinoma
C739|Thyroid_Gland|801|Carcinoma|8011/3|Malignant_Epithelioma
C739|Thyroid_Gland|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C739|Thyroid_Gland|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C739|Thyroid_Gland|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C739|Thyroid_Gland|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C739|Thyroid_Gland|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C739|Thyroid_Gland|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C739|Thyroid_Gland|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C739|Thyroid_Gland|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C739|Thyroid_Gland|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C739|Thyroid_Gland|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C739|Thyroid_Gland|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C739|Thyroid_Gland|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C739|Thyroid_Gland|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C739|Thyroid_Gland|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C739|Thyroid_Gland|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C739|Thyroid_Gland|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C739|Thyroid_Gland|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C739|Thyroid_Gland|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C739|Thyroid_Gland|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C739|Thyroid_Gland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C739|Thyroid_Gland|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C739|Thyroid_Gland|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C739|Thyroid_Gland|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C739|Thyroid_Gland|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C739|Thyroid_Gland|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C739|Thyroid_Gland|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C739|Thyroid_Gland|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C739|Thyroid_Gland|825|Bronchioloalveolar_Adenocarcinoma|8251/3|Bronchioloalveolar_Adenocarcinoma
C739|Thyroid_Gland|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C739|Thyroid_Gland|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C739|Thyroid_Gland|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C739|Thyroid_Gland|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C739|Thyroid_Gland|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C739|Thyroid_Gland|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C739|Thyroid_Gland|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C739|Thyroid_Gland|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C739|Thyroid_Gland|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C739|Thyroid_Gland|833|Follicular_Thyroid_Carcinoma|8330/3|Follicular_Thyroid_Carcinoma
C739|Thyroid_Gland|833|Follicular_Thyroid_Carcinoma|8331/3|Follicular_Thyroid_Carcinoma
C739|Thyroid_Gland|833|Follicular_Thyroid_Carcinoma|8332/3|Follicular_Thyroid_Carcinoma
C739|Thyroid_Gland|833|Follicular_Thyroid_Carcinoma|8333/3|Fetal_Adenocarcinoma
C739|Thyroid_Gland|833|Follicular_Thyroid_Carcinoma|8335/3|Follicular_Thyroid_Carcinoma
C739|Thyroid_Gland|833|Follicular_Thyroid_Carcinoma|8337/3|Poorly_Differentiated_Thyroid_Carcinoma
C739|Thyroid_Gland|833|Follicular_Thyroid_Carcinoma|8339/3|Follicular_Thyroid_Carcinoma
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8340/3|Papillary_Carcinoma__Follicular_Variant
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8341/3|Papillary_Microcarcinoma
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8342/3|Papillary_Carcinoma__Oxyphilic_Cell
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8343/2|Papillary_And_Follicular_Adenocarcinoma
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8343/3|Encapsulated_Papillary_Thyroid_Carcinoma
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8344/3|Papillary_Carcinoma__Columnar_Cell
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8345/3|Medullary_Carcinoma_With_Amyloid_Stroma
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8346/3|Mixed_Medullary_follicular_Carcinoma
C739|Thyroid_Gland|834|Papillary_And_Follicular_Adenocarcinoma|8347/3|Mixed_Medullary_papillary_Carcinoma
C739|Thyroid_Gland|835|Nonencapsulated_Sclerosing_Carcinoma|8350/3|Nonencapsulated_Sclerosing_Carcinoma
C739|Thyroid_Gland|845|Papillary_Cystadenocarcinoma|8450/3|Papillary_Cystadenocarcinoma
C739|Thyroid_Gland|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C739|Thyroid_Gland|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C739|Thyroid_Gland|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C739|Thyroid_Gland|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C739|Thyroid_Gland|898|Carcinosarcoma|8980/3|Carcinosarcoma
C739|Thyroid_Gland|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C739|Thyroid_Gland|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C739|Thyroid_Gland|959|Lymphoma|9590/3|Lymphoma
C739|Thyroid_Gland|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C739|Thyroid_Gland|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C739|Thyroid_Gland|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C739|Thyroid_Gland|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C739|Thyroid_Gland|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C739|Thyroid_Gland|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C739|Thyroid_Gland|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C739|Thyroid_Gland|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C739|Thyroid_Gland|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C739|Thyroid_Gland|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C739|Thyroid_Gland|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C739|Thyroid_Gland|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C739|Thyroid_Gland|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C739|Thyroid_Gland|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C739|Thyroid_Gland|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C739|Thyroid_Gland|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C739|Thyroid_Gland|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C739|Thyroid_Gland|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C739|Thyroid_Gland|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C739|Thyroid_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C739|Thyroid_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C739|Thyroid_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C739|Thyroid_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C739|Thyroid_Gland|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C739|Thyroid_Gland|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C739|Thyroid_Gland|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C739|Thyroid_Gland|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C739|Thyroid_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C739|Thyroid_Gland|970|T_Cell_Lymphoma|9701/3|Sezary_Syndrome
C739|Thyroid_Gland|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C739|Thyroid_Gland|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C739|Thyroid_Gland|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C739|Thyroid_Gland|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C739|Thyroid_Gland|971|Adult_Non_Hodgkin_Lymphoma|9715/3|Anaplastic_Large_Cell_Lymphoma
C739|Thyroid_Gland|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C739|Thyroid_Gland|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C739|Thyroid_Gland|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C739|Thyroid_Gland|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C739|Thyroid_Gland|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C739|Thyroid_Gland|973|Plasmacytoma|9731/3|Plasmacytoma
C739|Thyroid_Gland|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C739|Thyroid_Gland|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C739|Thyroid_Gland|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C739|Thyroid_Gland|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C739|Thyroid_Gland|974|Mast_Cell_Neoplasm|9740/3|Mast_Cell_Sarcoma
C739|Thyroid_Gland|974|Mast_Cell_Neoplasm|9741/3|Malignant_Mastocytosis
C739|Thyroid_Gland|974|Mast_Cell_Neoplasm|9749/3|Erdheim_Chester_Disease
C739|Thyroid_Gland|975|Neoplasm|9750/3|Malignant_Histiocytosis
C739|Thyroid_Gland|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C739|Thyroid_Gland|975|Neoplasm|9754/3|Adult_Langerhans_Cell_Histiocytosis
C739|Thyroid_Gland|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C739|Thyroid_Gland|975|Neoplasm|9756/3|Langerhans_Cell_Sarcoma
C739|Thyroid_Gland|975|Neoplasm|9757/3|Interdigitating_Dendritic_Cell_Sarcoma
C739|Thyroid_Gland|975|Neoplasm|9758/3|Follicular_Dendritic_Cell_Sarcoma
C739|Thyroid_Gland|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C739|Thyroid_Gland|976|Immunoproliferative_Disorder|9766/3|Lymphomatoid_Granulomatosis
C739|Thyroid_Gland|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C739|Thyroid_Gland|981|Neoplasm|9812/3|Lymphoma
C739|Thyroid_Gland|981|Neoplasm|9813/3|Lymphoma
C739|Thyroid_Gland|981|Neoplasm|9814/3|Lymphoma
C739|Thyroid_Gland|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C739|Thyroid_Gland|981|Neoplasm|9816/3|Hypodiploid_ALL
C739|Thyroid_Gland|981|Neoplasm|9817/3|Lymphoma
C739|Thyroid_Gland|981|Neoplasm|9818/3|Lymphoma
C739|Thyroid_Gland|981|Neoplasm|9819/3|Leukemia__B_Cell
C739|Thyroid_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C739|Thyroid_Gland|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C739|Thyroid_Gland|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C739|Thyroid_Gland|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C739|Thyroid_Gland|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C739|Thyroid_Gland|997|Neoplasm|9971/3|Polymorphic_PTLD
C739|Thyroid_Gland|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C740-C741,C749|Adrenal_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C740-C741,C749|Adrenal_Gland|800|Neoplasm|8001/3|Malignant_Cell
C740-C741,C749|Adrenal_Gland|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C740-C741,C749|Adrenal_Gland|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C740-C741,C749|Adrenal_Gland|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C740-C741,C749|Adrenal_Gland|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C740-C741,C749|Adrenal_Gland|801|Carcinoma|8010/2|In_Situ_Cancer
C740-C741,C749|Adrenal_Gland|801|Carcinoma|8010/3|Carcinoma
C740-C741,C749|Adrenal_Gland|801|Carcinoma|8011/3|Malignant_Epithelioma
C740-C741,C749|Adrenal_Gland|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C740-C741,C749|Adrenal_Gland|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C740-C741,C749|Adrenal_Gland|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C740-C741,C749|Adrenal_Gland|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C740-C741,C749|Adrenal_Gland|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C740-C741,C749|Adrenal_Gland|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C740-C741,C749|Adrenal_Gland|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C740-C741,C749|Adrenal_Gland|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C740-C741,C749|Adrenal_Gland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C740-C741,C749|Adrenal_Gland|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C740-C741,C749|Adrenal_Gland|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C740-C741,C749|Adrenal_Gland|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C740-C741,C749|Adrenal_Gland|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C740-C741,C749|Adrenal_Gland|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C740-C741,C749|Adrenal_Gland|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C740-C741,C749|Adrenal_Gland|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C740-C741,C749|Adrenal_Gland|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C740-C741,C749|Adrenal_Gland|837|Adrenocortical_Carcinoma|8370/3|Adrenocortical_Carcinoma
C740-C741,C749|Adrenal_Gland|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C740-C741,C749|Adrenal_Gland|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C740-C741,C749|Adrenal_Gland|870|Pheochromocytoma|8700/3|Pheochromocytoma
C740-C741,C749|Adrenal_Gland|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C740-C741,C749|Adrenal_Gland|906|Germ_Cell_Tumor|9064/3|Germinoma
C740-C741,C749|Adrenal_Gland|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C740-C741,C749|Adrenal_Gland|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C740-C741,C749|Adrenal_Gland|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C740-C741,C749|Adrenal_Gland|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C740-C741,C749|Adrenal_Gland|908|Teratoma|9080/3|Immature_Teratoma
C740-C741,C749|Adrenal_Gland|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C740-C741,C749|Adrenal_Gland|908|Teratoma|9082/3|Immature_Teratoma
C740-C741,C749|Adrenal_Gland|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C740-C741,C749|Adrenal_Gland|908|Teratoma|9084/3|Teratoma
C740-C741,C749|Adrenal_Gland|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C740-C741,C749|Adrenal_Gland|937|Chordoma|9370/3|Chordoma
C740-C741,C749|Adrenal_Gland|937|Chordoma|9371/3|Chondroid_Chordoma
C740-C741,C749|Adrenal_Gland|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C740-C741,C749|Adrenal_Gland|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C740-C741,C749|Adrenal_Gland|950|Neuroblastoma|9500/3|Neuroblastoma
C740-C741,C749|Adrenal_Gland|950|Neuroblastoma|9501/3|Medulloepithelioma
C740-C741,C749|Adrenal_Gland|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C740-C741,C749|Adrenal_Gland|950|Neuroblastoma|9503/3|Neuroepithelioma
C740-C741,C749|Adrenal_Gland|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C740-C741,C749|Adrenal_Gland|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C740-C741,C749|Adrenal_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C740-C741,C749|Adrenal_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C750|Parathyroid_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C750|Parathyroid_Gland|800|Neoplasm|8001/3|Malignant_Cell
C750|Parathyroid_Gland|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C750|Parathyroid_Gland|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C750|Parathyroid_Gland|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C750|Parathyroid_Gland|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C750|Parathyroid_Gland|801|Carcinoma|8010/2|In_Situ_Cancer
C750|Parathyroid_Gland|801|Carcinoma|8010/3|Carcinoma
C750|Parathyroid_Gland|801|Carcinoma|8011/3|Malignant_Epithelioma
C750|Parathyroid_Gland|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C750|Parathyroid_Gland|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C750|Parathyroid_Gland|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C750|Parathyroid_Gland|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C750|Parathyroid_Gland|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C750|Parathyroid_Gland|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C750|Parathyroid_Gland|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C750|Parathyroid_Gland|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C750|Parathyroid_Gland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C750|Parathyroid_Gland|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C750|Parathyroid_Gland|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C750|Parathyroid_Gland|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C750|Parathyroid_Gland|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C750|Parathyroid_Gland|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C750|Parathyroid_Gland|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C750|Parathyroid_Gland|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C750|Parathyroid_Gland|832|Granular_Cell_Carcinoma|8322/3|Water_Clear_Cell_Adenocarcinoma
C750|Parathyroid_Gland|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C750|Parathyroid_Gland|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C750|Parathyroid_Gland|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C750|Parathyroid_Gland|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C750|Parathyroid_Gland|906|Germ_Cell_Tumor|9064/3|Germinoma
C750|Parathyroid_Gland|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C750|Parathyroid_Gland|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C750|Parathyroid_Gland|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C750|Parathyroid_Gland|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C750|Parathyroid_Gland|908|Teratoma|9080/3|Immature_Teratoma
C750|Parathyroid_Gland|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C750|Parathyroid_Gland|908|Teratoma|9082/3|Immature_Teratoma
C750|Parathyroid_Gland|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C750|Parathyroid_Gland|908|Teratoma|9084/3|Teratoma
C750|Parathyroid_Gland|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C750|Parathyroid_Gland|937|Chordoma|9370/3|Chordoma
C750|Parathyroid_Gland|937|Chordoma|9371/3|Chondroid_Chordoma
C750|Parathyroid_Gland|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C750|Parathyroid_Gland|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C750|Parathyroid_Gland|950|Neuroblastoma|9500/3|Neuroblastoma
C750|Parathyroid_Gland|950|Neuroblastoma|9501/3|Medulloepithelioma
C750|Parathyroid_Gland|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C750|Parathyroid_Gland|950|Neuroblastoma|9503/3|Neuroepithelioma
C750|Parathyroid_Gland|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C750|Parathyroid_Gland|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C750|Parathyroid_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C750|Parathyroid_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C751|Pituitary_Gland|800|Neoplasm|8000/0|Benign_Neoplasm
C751|Pituitary_Gland|800|Neoplasm|8000/1|Neoplasm
C751|Pituitary_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C751|Pituitary_Gland|800|Neoplasm|8001/0|Tumor_Cells__Benign
C751|Pituitary_Gland|800|Neoplasm|8001/1|Neoplastic_Cell
C751|Pituitary_Gland|800|Neoplasm|8001/3|Malignant_Cell
C751|Pituitary_Gland|800|Neoplasm|8005/0|Clear_Cell_Neoplasm
C751|Pituitary_Gland|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C751|Pituitary_Gland|801|Carcinoma|8010/0|Benign_Epithelioma
C751|Pituitary_Gland|801|Carcinoma|8010/2|In_Situ_Cancer
C751|Pituitary_Gland|801|Carcinoma|8010/3|Carcinoma
C751|Pituitary_Gland|814|Adenocarcinoma|8140/0|Adenoma
C751|Pituitary_Gland|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C751|Pituitary_Gland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C751|Pituitary_Gland|814|Adenocarcinoma|8146/0|Salivary_Gland_Monomorphic_Adenoma
C751|Pituitary_Gland|826|Papillary_Adenocarcinoma|8260/0|Papillary_Adenoma
C751|Pituitary_Gland|827|Chromophobe_Renal_Cell_Carcinoma|8270/0|Pituitary_Gland_Chromophobe_Adenoma
C751|Pituitary_Gland|827|Chromophobe_Renal_Cell_Carcinoma|8270/3|Chromophobe_Renal_Cell_Carcinoma
C751|Pituitary_Gland|827|Chromophobe_Renal_Cell_Carcinoma|8271/0|Prolactinoma
C751|Pituitary_Gland|827|Chromophobe_Renal_Cell_Carcinoma|8272/0|Pituitary_Adenoma
C751|Pituitary_Gland|827|Chromophobe_Renal_Cell_Carcinoma|8272/3|Pituitary_Carcinoma
C751|Pituitary_Gland|827|Chromophobe_Renal_Cell_Carcinoma|8273/3|Blastoma
C751|Pituitary_Gland|828|Acidophil_Carcinoma|8280/0|Pituitary_Gland_Acidophil_Adenoma
C751|Pituitary_Gland|828|Acidophil_Carcinoma|8280/3|Acidophil_Carcinoma
C751|Pituitary_Gland|828|Acidophil_Carcinoma|8281/0|Mixed_Acidophil_basophil_Adenoma
C751|Pituitary_Gland|828|Acidophil_Carcinoma|8281/3|Mixed_Acidophil_basophil_Carcinoma
C751|Pituitary_Gland|829|Oxyphilic_Adenocarcinoma|8290/0|Oxyphilic_Adenoma
C751|Pituitary_Gland|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C751|Pituitary_Gland|830|Basophilic_Adenocarcinoma|8300/0|Pituitary_Gland_Basophil_Adenoma
C751|Pituitary_Gland|830|Basophilic_Adenocarcinoma|8300/3|Basophilic_Adenocarcinoma
C751|Pituitary_Gland|831|Clear_Cell_Adenocarcinoma|8310/0|Clear_Cell_Adenoma
C751|Pituitary_Gland|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C751|Pituitary_Gland|832|Granular_Cell_Carcinoma|8323/0|Mixed_Cell_Adenoma
C751|Pituitary_Gland|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C751|Pituitary_Gland|880|Sarcoma|8800/0|Benign_Soft_Tissue_Neoplasm
C751|Pituitary_Gland|880|Sarcoma|8800/3|Sarcoma
C751|Pituitary_Gland|885|Liposarcoma|8850/0|Lipoma
C751|Pituitary_Gland|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C751|Pituitary_Gland|906|Germ_Cell_Tumor|9064/3|Germinoma
C751|Pituitary_Gland|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C751|Pituitary_Gland|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C751|Pituitary_Gland|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C751|Pituitary_Gland|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C751|Pituitary_Gland|908|Teratoma|9080/0|Mature_Teratoma
C751|Pituitary_Gland|908|Teratoma|9080/1|Teratoma
C751|Pituitary_Gland|908|Teratoma|9080/3|Immature_Teratoma
C751|Pituitary_Gland|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C751|Pituitary_Gland|908|Teratoma|9082/3|Immature_Teratoma
C751|Pituitary_Gland|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C751|Pituitary_Gland|908|Teratoma|9084/3|Teratoma
C751|Pituitary_Gland|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C751|Pituitary_Gland|935|Craniopharyngioma|9350/1|Craniopharyngioma
C751|Pituitary_Gland|935|Craniopharyngioma|9351/1|Adamantinous_Craniopharyngioma
C751|Pituitary_Gland|935|Craniopharyngioma|9352/1|Papillary_Craniopharyngioma
C751|Pituitary_Gland|937|Chordoma|9370/3|Chordoma
C751|Pituitary_Gland|937|Chordoma|9371/3|Chondroid_Chordoma
C751|Pituitary_Gland|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C751|Pituitary_Gland|943|Astroblastoma|9432/1|Pituicytoma
C751|Pituitary_Gland|950|Neuroblastoma|9500/3|Neuroblastoma
C751|Pituitary_Gland|950|Neuroblastoma|9501/3|Medulloepithelioma
C751|Pituitary_Gland|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C751|Pituitary_Gland|950|Neuroblastoma|9503/3|Neuroepithelioma
C751|Pituitary_Gland|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C751|Pituitary_Gland|958|Granular_Cell_Tumor|9580/0|Granular_Cell_Tumor
C751|Pituitary_Gland|958|Granular_Cell_Tumor|9582/0|Granular_Cell_Tumor
C751|Pituitary_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C751|Pituitary_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C752|Craniopharyngeal_Duct|800|Neoplasm|8000/0|Benign_Neoplasm
C752|Craniopharyngeal_Duct|800|Neoplasm|8000/1|Neoplasm
C752|Craniopharyngeal_Duct|800|Neoplasm|8000/3|Malignant_Neoplasm
C752|Craniopharyngeal_Duct|800|Neoplasm|8001/0|Tumor_Cells__Benign
C752|Craniopharyngeal_Duct|800|Neoplasm|8001/1|Neoplastic_Cell
C752|Craniopharyngeal_Duct|800|Neoplasm|8001/3|Malignant_Cell
C752|Craniopharyngeal_Duct|800|Neoplasm|8005/0|Clear_Cell_Neoplasm
C752|Craniopharyngeal_Duct|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C752|Craniopharyngeal_Duct|801|Carcinoma|8010/0|Benign_Epithelioma
C752|Craniopharyngeal_Duct|801|Carcinoma|8010/2|In_Situ_Cancer
C752|Craniopharyngeal_Duct|801|Carcinoma|8010/3|Carcinoma
C752|Craniopharyngeal_Duct|814|Adenocarcinoma|8140/0|Adenoma
C752|Craniopharyngeal_Duct|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C752|Craniopharyngeal_Duct|814|Adenocarcinoma|8140/3|Adenocarcinoma
C752|Craniopharyngeal_Duct|814|Adenocarcinoma|8146/0|Salivary_Gland_Monomorphic_Adenoma
C752|Craniopharyngeal_Duct|826|Papillary_Adenocarcinoma|8260/0|Papillary_Adenoma
C752|Craniopharyngeal_Duct|827|Chromophobe_Renal_Cell_Carcinoma|8270/0|Pituitary_Gland_Chromophobe_Adenoma
C752|Craniopharyngeal_Duct|827|Chromophobe_Renal_Cell_Carcinoma|8270/3|Chromophobe_Renal_Cell_Carcinoma
C752|Craniopharyngeal_Duct|827|Chromophobe_Renal_Cell_Carcinoma|8271/0|Prolactinoma
C752|Craniopharyngeal_Duct|827|Chromophobe_Renal_Cell_Carcinoma|8272/0|Pituitary_Adenoma
C752|Craniopharyngeal_Duct|827|Chromophobe_Renal_Cell_Carcinoma|8272/3|Pituitary_Carcinoma
C752|Craniopharyngeal_Duct|828|Acidophil_Carcinoma|8280/0|Pituitary_Gland_Acidophil_Adenoma
C752|Craniopharyngeal_Duct|828|Acidophil_Carcinoma|8280/3|Acidophil_Carcinoma
C752|Craniopharyngeal_Duct|828|Acidophil_Carcinoma|8281/0|Mixed_Acidophil_basophil_Adenoma
C752|Craniopharyngeal_Duct|828|Acidophil_Carcinoma|8281/3|Mixed_Acidophil_basophil_Carcinoma
C752|Craniopharyngeal_Duct|829|Oxyphilic_Adenocarcinoma|8290/0|Oxyphilic_Adenoma
C752|Craniopharyngeal_Duct|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C752|Craniopharyngeal_Duct|830|Basophilic_Adenocarcinoma|8300/0|Pituitary_Gland_Basophil_Adenoma
C752|Craniopharyngeal_Duct|830|Basophilic_Adenocarcinoma|8300/3|Basophilic_Adenocarcinoma
C752|Craniopharyngeal_Duct|831|Clear_Cell_Adenocarcinoma|8310/0|Clear_Cell_Adenoma
C752|Craniopharyngeal_Duct|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C752|Craniopharyngeal_Duct|832|Granular_Cell_Carcinoma|8323/0|Mixed_Cell_Adenoma
C752|Craniopharyngeal_Duct|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C752|Craniopharyngeal_Duct|880|Sarcoma|8800/0|Benign_Soft_Tissue_Neoplasm
C752|Craniopharyngeal_Duct|880|Sarcoma|8800/3|Sarcoma
C752|Craniopharyngeal_Duct|885|Liposarcoma|8850/0|Lipoma
C752|Craniopharyngeal_Duct|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C752|Craniopharyngeal_Duct|906|Germ_Cell_Tumor|9064/3|Germinoma
C752|Craniopharyngeal_Duct|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C752|Craniopharyngeal_Duct|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C752|Craniopharyngeal_Duct|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C752|Craniopharyngeal_Duct|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C752|Craniopharyngeal_Duct|908|Teratoma|9080/0|Mature_Teratoma
C752|Craniopharyngeal_Duct|908|Teratoma|9080/1|Teratoma
C752|Craniopharyngeal_Duct|908|Teratoma|9080/3|Immature_Teratoma
C752|Craniopharyngeal_Duct|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C752|Craniopharyngeal_Duct|908|Teratoma|9082/3|Immature_Teratoma
C752|Craniopharyngeal_Duct|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C752|Craniopharyngeal_Duct|908|Teratoma|9084/3|Teratoma
C752|Craniopharyngeal_Duct|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C752|Craniopharyngeal_Duct|935|Craniopharyngioma|9350/1|Craniopharyngioma
C752|Craniopharyngeal_Duct|935|Craniopharyngioma|9351/1|Adamantinous_Craniopharyngioma
C752|Craniopharyngeal_Duct|935|Craniopharyngioma|9352/1|Papillary_Craniopharyngioma
C752|Craniopharyngeal_Duct|937|Chordoma|9370/3|Chordoma
C752|Craniopharyngeal_Duct|937|Chordoma|9371/3|Chondroid_Chordoma
C752|Craniopharyngeal_Duct|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C752|Craniopharyngeal_Duct|950|Neuroblastoma|9500/3|Neuroblastoma
C752|Craniopharyngeal_Duct|950|Neuroblastoma|9501/3|Medulloepithelioma
C752|Craniopharyngeal_Duct|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C752|Craniopharyngeal_Duct|950|Neuroblastoma|9503/3|Neuroepithelioma
C752|Craniopharyngeal_Duct|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C752|Craniopharyngeal_Duct|958|Granular_Cell_Tumor|9580/0|Granular_Cell_Tumor
C752|Craniopharyngeal_Duct|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C752|Craniopharyngeal_Duct|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C753|Pineal_Gland|800|Neoplasm|8000/0|Benign_Neoplasm
C753|Pineal_Gland|800|Neoplasm|8000/1|Neoplasm
C753|Pineal_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C753|Pineal_Gland|800|Neoplasm|8001/0|Tumor_Cells__Benign
C753|Pineal_Gland|800|Neoplasm|8001/1|Neoplastic_Cell
C753|Pineal_Gland|800|Neoplasm|8001/3|Malignant_Cell
C753|Pineal_Gland|801|Carcinoma|8010/0|Benign_Epithelioma
C753|Pineal_Gland|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C753|Pineal_Gland|906|Germ_Cell_Tumor|9064/3|Germinoma
C753|Pineal_Gland|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C753|Pineal_Gland|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C753|Pineal_Gland|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C753|Pineal_Gland|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C753|Pineal_Gland|908|Teratoma|9080/0|Mature_Teratoma
C753|Pineal_Gland|908|Teratoma|9080/3|Immature_Teratoma
C753|Pineal_Gland|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C753|Pineal_Gland|908|Teratoma|9082/3|Immature_Teratoma
C753|Pineal_Gland|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C753|Pineal_Gland|908|Teratoma|9084/0|Dermoid_Cyst
C753|Pineal_Gland|908|Teratoma|9084/3|Teratoma
C753|Pineal_Gland|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C753|Pineal_Gland|936|Neuroepithelioma__Peripheral|9360/1|Pineal_Gland_Neoplasm
C753|Pineal_Gland|936|Neuroepithelioma__Peripheral|9361/1|Pineocytoma
C753|Pineal_Gland|936|Neuroepithelioma__Peripheral|9362/3|Pineoblastoma
C753|Pineal_Gland|937|Chordoma|9370/3|Chordoma
C753|Pineal_Gland|937|Chordoma|9371/3|Chondroid_Chordoma
C753|Pineal_Gland|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C753|Pineal_Gland|939|Ependymoma|9395/3|Tumor_Of_The_Pineal_Region
C753|Pineal_Gland|947|Medulloblastoma|9473/3|Primitive_Neuroectodermal_Tumor
C753|Pineal_Gland|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C753|Pineal_Gland|949|Ganglioneuroblastoma|9492/0|Gangliocytoma
C753|Pineal_Gland|950|Neuroblastoma|9500/3|Neuroblastoma
C753|Pineal_Gland|950|Neuroblastoma|9501/3|Medulloepithelioma
C753|Pineal_Gland|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C753|Pineal_Gland|950|Neuroblastoma|9503/3|Neuroepithelioma
C753|Pineal_Gland|950|Neuroblastoma|9505/1|Ganglioglioma
C753|Pineal_Gland|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C753|Pineal_Gland|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C753|Pineal_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C753|Pineal_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C754-C755,C758-C759|Endocrine_Gland|800|Neoplasm|8000/3|Malignant_Neoplasm
C754-C755,C758-C759|Endocrine_Gland|800|Neoplasm|8001/3|Malignant_Cell
C754-C755,C758-C759|Endocrine_Gland|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C754-C755,C758-C759|Endocrine_Gland|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C754-C755,C758-C759|Endocrine_Gland|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C754-C755,C758-C759|Endocrine_Gland|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C754-C755,C758-C759|Endocrine_Gland|801|Carcinoma|8010/2|In_Situ_Cancer
C754-C755,C758-C759|Endocrine_Gland|801|Carcinoma|8010/3|Carcinoma
C754-C755,C758-C759|Endocrine_Gland|801|Carcinoma|8011/3|Malignant_Epithelioma
C754-C755,C758-C759|Endocrine_Gland|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C754-C755,C758-C759|Endocrine_Gland|814|Adenocarcinoma|8140/3|Adenocarcinoma
C754-C755,C758-C759|Endocrine_Gland|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C754-C755,C758-C759|Endocrine_Gland|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C754-C755,C758-C759|Endocrine_Gland|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C754-C755,C758-C759|Endocrine_Gland|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C754-C755,C758-C759|Endocrine_Gland|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C754-C755,C758-C759|Endocrine_Gland|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C754-C755,C758-C759|Endocrine_Gland|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C754-C755,C758-C759|Endocrine_Gland|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C754-C755,C758-C759|Endocrine_Gland|868|Paraganglioma|8681/3|Sympathetic_Paraganglioma
C754-C755,C758-C759|Endocrine_Gland|868|Paraganglioma|8682/3|Parasympathetic_Paraganglioma
C754-C755,C758-C759|Endocrine_Gland|869|Malignant_Extra_Adrenal_Paraganglioma|8690/3|Middle_Ear_Paraganglioma
C754-C755,C758-C759|Endocrine_Gland|869|Malignant_Extra_Adrenal_Paraganglioma|8691/3|Aorticopulmonary_Paraganglioma
C754-C755,C758-C759|Endocrine_Gland|869|Malignant_Extra_Adrenal_Paraganglioma|8692/3|Carotid_Body_Paraganglioma
C754-C755,C758-C759|Endocrine_Gland|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C754-C755,C758-C759|Endocrine_Gland|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C754-C755,C758-C759|Endocrine_Gland|906|Germ_Cell_Tumor|9064/3|Germinoma
C754-C755,C758-C759|Endocrine_Gland|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C754-C755,C758-C759|Endocrine_Gland|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C754-C755,C758-C759|Endocrine_Gland|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C754-C755,C758-C759|Endocrine_Gland|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C754-C755,C758-C759|Endocrine_Gland|908|Teratoma|9080/3|Immature_Teratoma
C754-C755,C758-C759|Endocrine_Gland|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C754-C755,C758-C759|Endocrine_Gland|908|Teratoma|9082/3|Immature_Teratoma
C754-C755,C758-C759|Endocrine_Gland|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C754-C755,C758-C759|Endocrine_Gland|908|Teratoma|9084/3|Teratoma
C754-C755,C758-C759|Endocrine_Gland|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C754-C755,C758-C759|Endocrine_Gland|937|Chordoma|9370/3|Chordoma
C754-C755,C758-C759|Endocrine_Gland|937|Chordoma|9371/3|Chondroid_Chordoma
C754-C755,C758-C759|Endocrine_Gland|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C754-C755,C758-C759|Endocrine_Gland|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C754-C755,C758-C759|Endocrine_Gland|950|Neuroblastoma|9500/3|Neuroblastoma
C754-C755,C758-C759|Endocrine_Gland|950|Neuroblastoma|9501/3|Medulloepithelioma
C754-C755,C758-C759|Endocrine_Gland|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C754-C755,C758-C759|Endocrine_Gland|950|Neuroblastoma|9503/3|Neuroepithelioma
C754-C755,C758-C759|Endocrine_Gland|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C754-C755,C758-C759|Endocrine_Gland|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C754-C755,C758-C759|Endocrine_Gland|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C754-C755,C758-C759|Endocrine_Gland|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C760-C768|Body_Region|800|Neoplasm|8000/3|Malignant_Neoplasm
C760-C768|Body_Region|800|Neoplasm|8001/3|Malignant_Cell
C760-C768|Body_Region|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C760-C768|Body_Region|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C760-C768|Body_Region|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C760-C768|Body_Region|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C760-C768|Body_Region|801|Carcinoma|8010/3|Carcinoma
C760-C768|Body_Region|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C760-C768|Body_Region|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C760-C768|Body_Region|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C760-C768|Body_Region|804|Non_Small_Cell_Carcinoma|8046/3|Non_Small_Cell_Carcinoma
C760-C768|Body_Region|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C760-C768|Body_Region|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C760-C768|Body_Region|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C760-C768|Body_Region|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C760-C768|Body_Region|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C760-C768|Body_Region|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C760-C768|Body_Region|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C760-C768|Body_Region|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C760-C768|Body_Region|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C760-C768|Body_Region|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C760-C768|Body_Region|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C760-C768|Body_Region|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C760-C768|Body_Region|814|Adenocarcinoma|8140/3|Adenocarcinoma
C760-C768|Body_Region|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C760-C768|Body_Region|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C760-C768|Body_Region|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C760-C768|Body_Region|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C760-C768|Body_Region|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C760-C768|Body_Region|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C760-C768|Body_Region|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C760-C768|Body_Region|845|Papillary_Cystadenocarcinoma|8450/3|Papillary_Cystadenocarcinoma
C760-C768|Body_Region|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C760-C768|Body_Region|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C760-C768|Body_Region|852|Intraductal_And_Lobular_Carcinoma|8525/3|Terminal_Duct_Adenocarcinoma
C760-C768|Body_Region|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C760-C768|Body_Region|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C760-C768|Body_Region|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C760-C768|Body_Region|950|Neuroblastoma|9500/3|Neuroblastoma
C760-C768|Body_Region|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C760-C768|Body_Region|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C770-C775,C778-C779|Lymph_Node|800|Neoplasm|8000/3|Malignant_Neoplasm
C770-C775,C778-C779|Lymph_Node|800|Neoplasm|8001/3|Malignant_Cell
C770-C775,C778-C779|Lymph_Node|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C770-C775,C778-C779|Lymph_Node|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C770-C775,C778-C779|Lymph_Node|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C770-C775,C778-C779|Lymph_Node|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C770-C775,C778-C779|Lymph_Node|959|Lymphoma|9590/3|Lymphoma
C770-C775,C778-C779|Lymph_Node|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C770-C775,C778-C779|Lymph_Node|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C770-C775,C778-C779|Lymph_Node|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C770-C775,C778-C779|Lymph_Node|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C770-C775,C778-C779|Lymph_Node|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C770-C775,C778-C779|Lymph_Node|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C770-C775,C778-C779|Lymph_Node|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C770-C775,C778-C779|Lymph_Node|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C770-C775,C778-C779|Lymph_Node|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C770-C775,C778-C779|Lymph_Node|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C770-C775,C778-C779|Lymph_Node|967|B_Cell_Lymphomas|9678/3|Primary_Effusion_Lymphoma
C770-C775,C778-C779|Lymph_Node|967|B_Cell_Lymphomas|9679/3|Mediastinal_Large_B_cell_Lymphoma
C770-C775,C778-C779|Lymph_Node|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C770-C775,C778-C779|Lymph_Node|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C770-C775,C778-C779|Lymph_Node|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C770-C775,C778-C779|Lymph_Node|968|Diffuse_Large_B_Cell_Lymphoma|9688/3|B_Cell_Non_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|968|Diffuse_Large_B_Cell_Lymphoma|9689/3|Mucosa_associated_Lymphoma
C770-C775,C778-C779|Lymph_Node|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C770-C775,C778-C779|Lymph_Node|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C770-C775,C778-C779|Lymph_Node|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C770-C775,C778-C779|Lymph_Node|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C770-C775,C778-C779|Lymph_Node|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C770-C775,C778-C779|Lymph_Node|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C770-C775,C778-C779|Lymph_Node|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C770-C775,C778-C779|Lymph_Node|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C770-C775,C778-C779|Lymph_Node|971|Adult_Non_Hodgkin_Lymphoma|9712/3|Angioendotheliomatosis
C770-C775,C778-C779|Lymph_Node|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C770-C775,C778-C779|Lymph_Node|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C770-C775,C778-C779|Lymph_Node|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C770-C775,C778-C779|Lymph_Node|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C770-C775,C778-C779|Lymph_Node|972|Lymphoblastic_Lymphoma|9724/3|Lymphoproliferative_Disorder
C770-C775,C778-C779|Lymph_Node|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C770-C775,C778-C779|Lymph_Node|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C770-C775,C778-C779|Lymph_Node|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C770-C775,C778-C779|Lymph_Node|973|Plasmacytoma|9735/3|Plasmablastic_Lymphoma
C770-C775,C778-C779|Lymph_Node|973|Plasmacytoma|9737/3|B_Cell_Non_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|973|Plasmacytoma|9738/3|B_Cell_Non_Hodgkin_Lymphoma
C770-C775,C778-C779|Lymph_Node|975|Neoplasm|9751/3|Adult_Langerhans_Cell_Histiocytosis
C770-C775,C778-C779|Lymph_Node|975|Neoplasm|9755/3|Histiocytic_Sarcoma
C770-C775,C778-C779|Lymph_Node|975|Neoplasm|9759/3|Fibroblastic_Reticular_Cell_Tumor
C770-C775,C778-C779|Lymph_Node|976|Immunoproliferative_Disorder|9761/3|Waldenstrom_Macroglobulinemia
C770-C775,C778-C779|Lymph_Node|976|Immunoproliferative_Disorder|9762/3|Heavy_Chain_Disease
C770-C775,C778-C779|Lymph_Node|981|Neoplasm|9811/3|B_Lymphoblastic_Leukemia_Lymphoma
C770-C775,C778-C779|Lymph_Node|981|Neoplasm|9812/3|Lymphoma
C770-C775,C778-C779|Lymph_Node|981|Neoplasm|9813/3|Lymphoma
C770-C775,C778-C779|Lymph_Node|981|Neoplasm|9814/3|Lymphoma
C770-C775,C778-C779|Lymph_Node|981|Neoplasm|9815/3|B_Lymphoblastic_Leukemia_Lymphoma
C770-C775,C778-C779|Lymph_Node|981|Neoplasm|9816/3|Hypodiploid_ALL
C770-C775,C778-C779|Lymph_Node|981|Neoplasm|9817/3|Lymphoma
C770-C775,C778-C779|Lymph_Node|981|Neoplasm|9818/3|Lymphoma
C770-C775,C778-C779|Lymph_Node|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
C770-C775,C778-C779|Lymph_Node|983|Leukemia|9831/3|Leukemia__Large_Granular_Lymphocytic
C770-C775,C778-C779|Lymph_Node|983|Leukemia|9837/3|T_Lymphoblastic_Leukemia_Lymphoma
C770-C775,C778-C779|Lymph_Node|996|Myeloproliferative_Neoplasm|9965/3|Neoplasm
C770-C775,C778-C779|Lymph_Node|996|Myeloproliferative_Neoplasm|9967/3|Lymphocytic_Neoplasm
C770-C775,C778-C779|Lymph_Node|997|Neoplasm|9971/3|Polymorphic_PTLD
C770-C775,C778-C779|Lymph_Node|997|Neoplasm|9975/3|Myeloproliferative_Neoplasm
C809|Body_Region|800|Neoplasm|8000/3|Malignant_Neoplasm
C809|Body_Region|800|Neoplasm|8001/3|Malignant_Cell
C809|Body_Region|800|Neoplasm|8002/3|Malignant_Tumor__Small_Cell_Type
C809|Body_Region|800|Neoplasm|8003/3|Malignant_Giant_Cell_Neoplasm
C809|Body_Region|800|Neoplasm|8004/3|Malignant_Spindle_Cell_Neoplasm
C809|Body_Region|800|Neoplasm|8005/3|Malignant_Tumor__Clear_Cell_Type
C809|Body_Region|801|Carcinoma|8010/2|In_Situ_Cancer
C809|Body_Region|801|Carcinoma|8010/3|Carcinoma
C809|Body_Region|801|Carcinoma|8011/3|Malignant_Epithelioma
C809|Body_Region|801|Carcinoma|8012/3|Large_Cell_Carcinoma
C809|Body_Region|801|Carcinoma|8013/3|Large_Cell_Neuroendocrine_Carcinoma
C809|Body_Region|801|Carcinoma|8014/3|Large_Cell_Carcinoma
C809|Body_Region|801|Carcinoma|8015/3|Glassy_Cell_Carcinoma
C809|Body_Region|802|Carcinoma|8020/3|Undifferentiated_Carcinoma
C809|Body_Region|802|Carcinoma|8021/3|Undifferentiated_Carcinoma
C809|Body_Region|802|Carcinoma|8022/3|Pleomorphic_Carcinoma
C809|Body_Region|803|Sarcomatoid_Carcinoma|8030/3|Giant_Cell_And_Spindle_Cell_Carcinoma
C809|Body_Region|803|Sarcomatoid_Carcinoma|8031/3|Giant_Cell_Carcinoma
C809|Body_Region|803|Sarcomatoid_Carcinoma|8032/3|Sarcomatoid_Carcinoma
C809|Body_Region|803|Sarcomatoid_Carcinoma|8033/3|Sarcomatoid_Carcinoma
C809|Body_Region|803|Sarcomatoid_Carcinoma|8034/3|Polygonal_Cell_Carcinoma
C809|Body_Region|803|Sarcomatoid_Carcinoma|8035/3|Carcinoma
C809|Body_Region|804|Small_Cell_Carcinoma|8041/3|Small_Cell_Carcinoma
C809|Body_Region|804|Small_Cell_Carcinoma|8043/3|Small_Cell_Carcinoma__Fusiform_Cell
C809|Body_Region|805|Papillary_Carcinoma|8050/2|Papillary_Carcinoma_In_Situ
C809|Body_Region|805|Papillary_Carcinoma|8050/3|Papillary_Carcinoma
C809|Body_Region|805|Papillary_Carcinoma|8051/3|Verrucous_Carcinoma
C809|Body_Region|805|Papillary_Carcinoma|8052/2|Papillary_Squamous_Cell_Carcinoma
C809|Body_Region|805|Papillary_Carcinoma|8052/3|Papillary_Squamous_Cell_Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8070/2|Stage_0_Squamous_Cell_Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8070/3|Squamous_Cell_Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8071/3|Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8072/3|Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8073/3|Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8074/3|Sarcomatoid_Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8075/3|Pseudoglandular_Squamous_Cell_Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8076/2|Stage_0_Squamous_Cell_Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8076/3|Carcinoma
C809|Body_Region|807|Squamous_Cell_Carcinoma|8078/3|Squamous_Cell_Carcinoma
C809|Body_Region|808|Lymphoepithelial_Carcinoma|8082/3|Lymphoepithelial_Carcinoma
C809|Body_Region|808|Lymphoepithelial_Carcinoma|8083/3|Basaloid_Squamous_Cell_Carcinoma
C809|Body_Region|808|Lymphoepithelial_Carcinoma|8084/3|Squamous_Cell_Carcinoma
C809|Body_Region|812|Transitional_Cell_Carcinoma|8120/2|Stage_0_Transitional_Cell_Carcinoma
C809|Body_Region|812|Transitional_Cell_Carcinoma|8120/3|Transitional_Cell_Carcinoma
C809|Body_Region|812|Transitional_Cell_Carcinoma|8121/3|Schneiderian_Carcinoma
C809|Body_Region|812|Transitional_Cell_Carcinoma|8122/3|Sarcomatoid_Carcinoma
C809|Body_Region|812|Transitional_Cell_Carcinoma|8123/3|Basaloid_Carcinoma
C809|Body_Region|812|Transitional_Cell_Carcinoma|8124/3|Anal_Canal_Cloacogenic_Carcinoma
C809|Body_Region|813|Carcinoma|8130/2|Carcinoma
C809|Body_Region|813|Carcinoma|8130/3|Carcinoma
C809|Body_Region|813|Carcinoma|8131/3|Transitional_Cell_Carcinoma
C809|Body_Region|814|Adenocarcinoma|8140/2|Adenocarcinoma_In_Situ
C809|Body_Region|814|Adenocarcinoma|8140/3|Adenocarcinoma
C809|Body_Region|814|Adenocarcinoma|8141/3|Scirrhous_Adenocarcinoma
C809|Body_Region|814|Adenocarcinoma|8143/3|Superficial_Spreading_Adenocarcinoma
C809|Body_Region|814|Adenocarcinoma|8147/3|Adenocarcinoma__Basal_Cell
C809|Body_Region|815|Endocrine_Gland_Neoplasms|8152/3|Malignant_Pancreatic_Glucagonoma
C809|Body_Region|815|Endocrine_Gland_Neoplasms|8153/3|Malignant_Gastrinoma
C809|Body_Region|815|Endocrine_Gland_Neoplasms|8156/3|Malignant_Somatostatinoma
C809|Body_Region|815|Endocrine_Gland_Neoplasms|8157/3|Malignant_Enteroglucagonoma
C809|Body_Region|819|Trabecular_Adenocarcinoma|8190/3|Trabecular_Adenocarcinoma
C809|Body_Region|820|Cribriform_Carcinoma|8200/3|Adenoid_Cystic_Carcinoma
C809|Body_Region|820|Cribriform_Carcinoma|8201/2|Cribriform_Carcinoma_In_Situ
C809|Body_Region|820|Cribriform_Carcinoma|8201/3|Cribriform_Carcinoma
C809|Body_Region|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/2|Adenocarcinoma_In_Situ
C809|Body_Region|821|Adenocarcinoma_In_Adenomatous_Polyp|8210/3|Adenocarcinoma_In_Adenomatous_Polyp
C809|Body_Region|821|Adenocarcinoma_In_Adenomatous_Polyp|8211/3|Tubular_Adenocarcinoma
C809|Body_Region|823|Solid_Carcinoma|8230/2|In_Situ_Cancer
C809|Body_Region|823|Solid_Carcinoma|8230/3|Solid_Carcinoma
C809|Body_Region|823|Solid_Carcinoma|8231/3|Carcinoma_Simplex
C809|Body_Region|824|Atypical_Carcinoid_Tumor|8240/3|Atypical_Carcinoid_Tumor
C809|Body_Region|824|Atypical_Carcinoid_Tumor|8241/3|EC_Cell_Carcinoid
C809|Body_Region|824|Atypical_Carcinoid_Tumor|8242/3|Malignant_Neoplasm
C809|Body_Region|824|Atypical_Carcinoid_Tumor|8243/3|Goblet_Cell_Carcinoid
C809|Body_Region|824|Atypical_Carcinoid_Tumor|8244/3|Adenocarcinoid_Tumor
C809|Body_Region|824|Atypical_Carcinoid_Tumor|8245/3|Adenocarcinoid_Tumor
C809|Body_Region|824|Atypical_Carcinoid_Tumor|8246/3|Carcinoma__Neuroendocrine
C809|Body_Region|824|Atypical_Carcinoid_Tumor|8249/3|Atypical_Carcinoid_Tumor
C809|Body_Region|825|Bronchioloalveolar_Adenocarcinoma|8251/3|Bronchioloalveolar_Adenocarcinoma
C809|Body_Region|825|Bronchioloalveolar_Adenocarcinoma|8255/3|Adenocarcinoma_With_Mixed_Subtypes
C809|Body_Region|826|Papillary_Adenocarcinoma|8260/3|Papillary_Adenocarcinoma
C809|Body_Region|826|Papillary_Adenocarcinoma|8261/2|Adenocarcinoma_In_Situ
C809|Body_Region|826|Papillary_Adenocarcinoma|8261/3|Adenocarcinoma_In_Villous_Adenoma
C809|Body_Region|826|Papillary_Adenocarcinoma|8262/3|Villous_Adenocarcinoma
C809|Body_Region|826|Papillary_Adenocarcinoma|8263/2|Adenocarcinoma_In_Situ
C809|Body_Region|826|Papillary_Adenocarcinoma|8263/3|Adenocarcinoma_In_Tubulovillous_Adenoma
C809|Body_Region|829|Oxyphilic_Adenocarcinoma|8290/3|Oxyphilic_Adenocarcinoma
C809|Body_Region|831|Clear_Cell_Adenocarcinoma|8310/3|Clear_Cell_Adenocarcinoma
C809|Body_Region|832|Granular_Cell_Carcinoma|8320/3|Granular_Cell_Carcinoma
C809|Body_Region|832|Granular_Cell_Carcinoma|8323/3|Mixed_Cell_Adenocarcinoma
C809|Body_Region|838|Carcinoma__Endometrioid|8380/3|Carcinoma__Endometrioid
C809|Body_Region|840|Sweat_Gland_Adenocarcinoma|8401/3|Apocrine_Adenocarcinoma
C809|Body_Region|843|Mucoepidermoid_Carcinoma|8430/3|Mucoepidermoid_Carcinoma
C809|Body_Region|844|Cystadenocarcinoma|8440/3|Cystadenocarcinoma
C809|Body_Region|848|Mucinous_Adenocarcinoma|8480/3|Mucinous_Adenocarcinoma
C809|Body_Region|848|Mucinous_Adenocarcinoma|8481/3|Mucin_Producing_Adenocarcinoma
C809|Body_Region|849|Signet_Ring_Cell_Carcinoma|8490/3|Signet_Ring_Cell_Carcinoma
C809|Body_Region|851|Medullary_Carcinoma|8510/3|Medullary_Carcinoma
C809|Body_Region|852|Intraductal_And_Lobular_Carcinoma|8521/3|Invasive_Ductal_Breast_Carcinoma
C809|Body_Region|854|Paget_Disease_Extramammary|8542/3|Paget_Disease_Extramammary
C809|Body_Region|855|Acinar_Cell_Carcinoma|8550/3|Acinar_Cell_Carcinoma
C809|Body_Region|855|Acinar_Cell_Carcinoma|8551/3|Acinar_Cell_Cystadenocarcinoma
C809|Body_Region|856|Adenosquamous_Carcinoma|8560/3|Adenosquamous_Carcinoma
C809|Body_Region|856|Adenosquamous_Carcinoma|8562/3|Epithelial_Myoepithelial_Carcinoma
C809|Body_Region|857|Adenocarcinoma_With_Metaplasia|8570/3|Adenocarcinoma_With_Squamous_Metaplasia
C809|Body_Region|857|Adenocarcinoma_With_Metaplasia|8571/3|Adenocarcinoma
C809|Body_Region|857|Adenocarcinoma_With_Metaplasia|8572/3|Adenocarcinoma
C809|Body_Region|857|Adenocarcinoma_With_Metaplasia|8573/3|Adenocarcinoma_With_Apocrine_Metaplasia
C809|Body_Region|857|Adenocarcinoma_With_Metaplasia|8574/3|Adenocarcinoma
C809|Body_Region|857|Adenocarcinoma_With_Metaplasia|8575/3|Metaplastic_Carcinoma
C809|Body_Region|863|Neoplasm|8630/3|Malignant_Sertoli_Cell_Tumor
C809|Body_Region|865|Malignant_Leydig_Cell_Tumor|8650/3|Malignant_Leydig_Cell_Tumor
C809|Body_Region|868|Paraganglioma|8680/3|Malignant_Paraganglioma
C809|Body_Region|869|Malignant_Extra_Adrenal_Paraganglioma|8693/3|Malignant_Extra_Adrenal_Paraganglioma
C809|Body_Region|871|Malignant_Glomus_Tumor|8710/3|Malignant_Glomus_Tumor
C809|Body_Region|880|Sarcoma|8800/3|Sarcoma
C809|Body_Region|880|Sarcoma|8801/3|Spindle_Cell_Sarcoma
C809|Body_Region|880|Sarcoma|8802/3|Giant_Cell_Sarcoma
C809|Body_Region|880|Sarcoma|8803/3|Small_Cell_Sarcoma
C809|Body_Region|880|Sarcoma|8804/3|Sarcoma__Epithelioid
C809|Body_Region|880|Sarcoma|8805/3|Undifferentiated_Sarcoma
C809|Body_Region|880|Sarcoma|8806/3|Desmoplastic_Small_Round_Cell_Tumor
C809|Body_Region|881|Fibromatous_Neoplasm|8810/3|Fibrosarcoma
C809|Body_Region|881|Fibromatous_Neoplasm|8811/3|Myxofibrosarcoma
C809|Body_Region|881|Fibromatous_Neoplasm|8813/3|Fascial_Fibrosarcoma
C809|Body_Region|881|Fibromatous_Neoplasm|8814/3|Infantile_Fibrosarcoma
C809|Body_Region|881|Fibromatous_Neoplasm|8815/3|Malignant_Solitary_Fibrous_Tumor
C809|Body_Region|882|Sarcoma|8825/3|Sarcoma
C809|Body_Region|883|Benign_Fibrous_Histiocytoma|8830/3|Malignant_Fibrous_Histiocytoma
C809|Body_Region|884|Myxosarcoma|8840/3|Myxosarcoma
C809|Body_Region|885|Liposarcoma|8850/3|Liposarcoma
C809|Body_Region|885|Liposarcoma|8851/3|Well_Differentiated_Liposarcoma
C809|Body_Region|885|Liposarcoma|8852/3|Liposarcoma__Myxoid
C809|Body_Region|885|Liposarcoma|8853/3|Round_Cell_Liposarcoma
C809|Body_Region|885|Liposarcoma|8854/3|Pleomorphic_Liposarcoma
C809|Body_Region|885|Liposarcoma|8855/3|Liposarcoma
C809|Body_Region|885|Liposarcoma|8857/3|Fibroblastic_Liposarcoma
C809|Body_Region|885|Liposarcoma|8858/3|Dedifferentiated_Liposarcoma
C809|Body_Region|889|Myomatous_Neoplasm|8890/3|Leiomyosarcoma
C809|Body_Region|889|Myomatous_Neoplasm|8891/3|Epithelioid_Leiomyosarcoma
C809|Body_Region|889|Myomatous_Neoplasm|8894/3|Angiomyosarcoma
C809|Body_Region|889|Myomatous_Neoplasm|8895/3|Myosarcoma
C809|Body_Region|889|Myomatous_Neoplasm|8896/3|Myxoid_Leiomyosarcoma
C809|Body_Region|890|Rhabdomyosarcoma|8900/3|Rhabdomyosarcoma
C809|Body_Region|890|Rhabdomyosarcoma|8901/3|Pleomorphic_Rhabdomyosarcoma
C809|Body_Region|890|Rhabdomyosarcoma|8902/3|Mixed_Type_Rhabdomyosarcoma
C809|Body_Region|891|Embryonal_Rhabdomyosarcoma|8910/3|Embryonal_Rhabdomyosarcoma
C809|Body_Region|891|Embryonal_Rhabdomyosarcoma|8912/3|Spindle_Cell_Rhabdomyosarcoma
C809|Body_Region|892|Alveolar_Rhabdomyosarcoma|8920/3|Alveolar_Rhabdomyosarcoma
C809|Body_Region|892|Alveolar_Rhabdomyosarcoma|8921/3|Rhabdomyosarcoma
C809|Body_Region|893|Stromal_Sarcoma|8934/3|Carcinofibroma
C809|Body_Region|893|Stromal_Sarcoma|8935/3|Stromal_Sarcoma
C809|Body_Region|894|Malignant_Mixed_Tumor|8940/3|Malignant_Mixed_Tumor
C809|Body_Region|894|Malignant_Mixed_Tumor|8941/3|Carcinoma_Ex_Pleomorphic_Adenoma
C809|Body_Region|895|Mixed_Tumor__Mullerian|8950/3|Mixed_Tumor__Mullerian
C809|Body_Region|895|Mixed_Tumor__Mullerian|8951/3|Mesodermal_Mixed_Tumor
C809|Body_Region|898|Carcinosarcoma|8980/3|Carcinosarcoma
C809|Body_Region|898|Carcinosarcoma|8981/3|Carcinosarcoma__Embryonal
C809|Body_Region|898|Carcinosarcoma|8982/3|Malignant_Myoepithelioma
C809|Body_Region|899|Malignant_Mesenchymoma|8990/3|Malignant_Mesenchymoma
C809|Body_Region|899|Malignant_Mesenchymoma|8991/3|Undifferentiated__Embryonal__Sarcoma
C809|Body_Region|904|Synovial_Sarcoma|9040/3|Synovial_Sarcoma
C809|Body_Region|904|Synovial_Sarcoma|9041/3|Spindle_Cell_Synovial_Sarcoma
C809|Body_Region|904|Synovial_Sarcoma|9042/3|Epithelial_Synovial_Sarcoma
C809|Body_Region|904|Synovial_Sarcoma|9043/3|Biphasic_Synovial_Sarcoma
C809|Body_Region|904|Synovial_Sarcoma|9044/3|Clear_Cell_Sarcoma_Of_Soft_Tissue_C0206651
C809|Body_Region|906|Germ_Cell_Tumor|9060/3|Dysgerminoma
C809|Body_Region|906|Germ_Cell_Tumor|9064/3|Germinoma
C809|Body_Region|906|Germ_Cell_Tumor|9065/3|Nongerminomatous_Germ_Cell_Tumor_C1266158
C809|Body_Region|907|Embryonal_Carcinoma|9070/3|Embryonal_Carcinoma
C809|Body_Region|907|Embryonal_Carcinoma|9071/3|Yolk_Sac_Tumor
C809|Body_Region|907|Embryonal_Carcinoma|9072/3|Polyembryoma
C809|Body_Region|908|Teratoma|9080/3|Immature_Teratoma
C809|Body_Region|908|Teratoma|9081/3|Mixed_Embryonal_Carcinoma_And_Teratoma
C809|Body_Region|908|Teratoma|9082/3|Immature_Teratoma
C809|Body_Region|908|Teratoma|9083/3|Intermediate_Immature_Teratoma
C809|Body_Region|908|Teratoma|9084/3|Teratoma
C809|Body_Region|908|Teratoma|9085/3|Mixed_Germ_Cell_Tumor
C809|Body_Region|910|Choriocarcinoma|9100/3|Choriocarcinoma
C809|Body_Region|910|Choriocarcinoma|9101/3|Choriocarcinoma
C809|Body_Region|910|Choriocarcinoma|9102/3|Malignant_Trophoblastic_Teratoma
C809|Body_Region|910|Choriocarcinoma|9105/3|Epithelioid_Trophoblastic_Tumor
C809|Body_Region|911|Mesonephroma|9110/3|Mesonephroma
C809|Body_Region|912|Neoplasms__Vascular_Tissue|9120/3|Hemangiosarcoma
C809|Body_Region|913|Hemangioendothelioma|9130/3|Hemangiosarcoma
C809|Body_Region|913|Hemangioendothelioma|9133/3|Epithelioid_Hemangioendothelioma
C809|Body_Region|914|Kaposi_Sarcoma|9140/3|Kaposi_Sarcoma
C809|Body_Region|915|Hemangiopericytoma|9150/3|Malignant_Hemangiopericytoma
C809|Body_Region|917|Lymphangiosarcoma|9170/3|Lymphangiosarcoma
C809|Body_Region|931|Malignant_Ameloblastoma|9310/3|Malignant_Ameloblastoma
C809|Body_Region|937|Chordoma|9370/3|Chordoma
C809|Body_Region|937|Chordoma|9371/3|Chondroid_Chordoma
C809|Body_Region|937|Chordoma|9372/3|Dedifferentiated_Chordoma
C809|Body_Region|949|Ganglioneuroblastoma|9490/3|Ganglioneuroblastoma
C809|Body_Region|950|Neuroblastoma|9500/3|Neuroblastoma
C809|Body_Region|950|Neuroblastoma|9501/3|Medulloepithelioma
C809|Body_Region|950|Neuroblastoma|9502/3|Teratoid_Medulloepithelioma
C809|Body_Region|950|Neuroblastoma|9503/3|Neuroepithelioma
C809|Body_Region|950|Neuroblastoma|9504/3|Polar_Spongioblastoma
C809|Body_Region|950|Neuroblastoma|9505/3|Anaplastic_Ganglioglioma
C809|Body_Region|952|Neoplasm|9520/3|Neoplasm
C809|Body_Region|954|Malignant_Peripheral_Nerve_Sheath_Tumor|9540/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C809|Body_Region|956|Schwannoma|9560/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C809|Body_Region|956|Schwannoma|9561/3|Malignant_Peripheral_Nerve_Sheath_Tumor
C809|Body_Region|957|Perineurioma|9571/3|Malignant_Perineurioma
C809|Body_Region|958|Granular_Cell_Tumor|9580/3|Malignant_Granular_Cell_Tumor
C809|Body_Region|958|Granular_Cell_Tumor|9581/3|Alveolar_Soft_Part_Sarcoma
C809|Body_Region|959|Lymphoma|9590/3|Lymphoma
C809|Body_Region|959|Lymphoma|9591/3|Adult_Non_Hodgkin_Lymphoma
C809|Body_Region|959|Lymphoma|9596/3|Adult_Non_Hodgkin_Lymphoma
C809|Body_Region|965|Adult_Hodgkin_Lymphoma|9650/3|Adult_Hodgkin_Lymphoma
C809|Body_Region|965|Adult_Hodgkin_Lymphoma|9651/3|Hodgkin_Lymphoma__Lymphocyte_rich
C809|Body_Region|965|Adult_Hodgkin_Lymphoma|9652/3|Mixed_Cellularity_Hodgkin_Lymphoma
C809|Body_Region|965|Adult_Hodgkin_Lymphoma|9653/3|Chronic_Lymphocytic_Leukemia
C809|Body_Region|965|Adult_Hodgkin_Lymphoma|9654/3|Hodgkin_Lymphoma__Lymphocyte_Depletion
C809|Body_Region|965|Adult_Hodgkin_Lymphoma|9655/3|Adult_Hodgkin_Lymphoma
C809|Body_Region|965|Adult_Hodgkin_Lymphoma|9659/3|Childhood_NLPHD
C809|Body_Region|966|Adult_Hodgkin_Lymphoma|9661/3|Hodgkin_s_Granuloma
C809|Body_Region|966|Adult_Hodgkin_Lymphoma|9662/3|Adult_Hodgkin_Lymphoma
C809|Body_Region|966|Adult_Hodgkin_Lymphoma|9663/3|Hodgkin_s_Nodular_Sclerosis
C809|Body_Region|966|Adult_Hodgkin_Lymphoma|9664/3|Adult_Hodgkin_Lymphoma
C809|Body_Region|966|Adult_Hodgkin_Lymphoma|9665/3|Adult_Hodgkin_Lymphoma
C809|Body_Region|966|Adult_Hodgkin_Lymphoma|9667/3|Adult_Hodgkin_Lymphoma
C809|Body_Region|967|B_Cell_Lymphomas|9670/3|Small_Lymphocytic_Lymphoma
C809|Body_Region|967|B_Cell_Lymphomas|9671/3|Lymphoplasmacytic_Lymphoma
C809|Body_Region|967|B_Cell_Lymphomas|9673/3|Mantle_Cell_Lymphoma
C809|Body_Region|967|B_Cell_Lymphomas|9675/3|Diffuse_Malignant_Lymphoma
C809|Body_Region|967|B_Cell_Lymphomas|9678/3|Primary_Effusion_Lymphoma
C809|Body_Region|967|B_Cell_Lymphomas|9679/3|Mediastinal_Large_B_cell_Lymphoma
C809|Body_Region|968|Diffuse_Large_B_Cell_Lymphoma|9680/3|Diffuse_Large_B_Cell_Lymphoma
C809|Body_Region|968|Diffuse_Large_B_Cell_Lymphoma|9684/3|Immunoblastic_Lymphoma
C809|Body_Region|968|Diffuse_Large_B_Cell_Lymphoma|9687/3|Burkitt_Lymphoma
C809|Body_Region|968|Diffuse_Large_B_Cell_Lymphoma|9689/3|Mucosa_associated_Lymphoma
C809|Body_Region|969|Follicular_Adenoma|9690/3|Lymphoma__Follicular
C809|Body_Region|969|Follicular_Adenoma|9691/3|Grade_2_Follicular_Lymphoma
C809|Body_Region|969|Follicular_Adenoma|9695/3|Follicular_Lymphoma__Grade_1
C809|Body_Region|969|Follicular_Adenoma|9698/3|Lymphoma__Follicular__Grade_3
C809|Body_Region|969|Follicular_Adenoma|9699/3|Mucosa_associated_Lymphoma
C809|Body_Region|970|T_Cell_Lymphoma|9702/3|Peripheral_T_Cell_Lymphoma
C809|Body_Region|970|T_Cell_Lymphoma|9705/3|Angioimmunoblastic_Lymphadenopathy
C809|Body_Region|970|T_Cell_Lymphoma|9708/3|T_Cell_Lymphoma
C809|Body_Region|971|Adult_Non_Hodgkin_Lymphoma|9714/3|Anaplastic_Large_Cell_Lymphoma
C809|Body_Region|971|Adult_Non_Hodgkin_Lymphoma|9716/3|Lymphoma
C809|Body_Region|971|Adult_Non_Hodgkin_Lymphoma|9717/3|Intestinal_T_Cell_Lymphoma__NOS
C809|Body_Region|971|Adult_Non_Hodgkin_Lymphoma|9719/3|T_Cell_Lymphoma
C809|Body_Region|972|Lymphoblastic_Lymphoma|9727/3|Lymphoblastic_Lymphoma
C809|Body_Region|972|Lymphoblastic_Lymphoma|9728/3|Lymphoblastic_Lymphoma
C809|Body_Region|972|Lymphoblastic_Lymphoma|9729/3|Lymphoblastic_Lymphoma
C809|Body_Region|973|Plasmacytoma|9731/3|Plasmacytoma
C809|Body_Region|973|Plasmacytoma|9732/3|Plasma_Cell_Myeloma
C809|Body_Region|973|Plasmacytoma|9734/3|Extramedullary_Plasmacytoma
C809|Body_Region|982|Lymphoid_Leukemia|9823/3|Chronic_Lymphocytic_Leukemia
