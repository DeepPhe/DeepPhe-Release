Alpha Or Number Description Colon||^[ \t]*(?<Index>[A-Z0-9])[\).:][ \t]+(?<Subject>[^:\r\n]+):[ \t]*\r?\n
Alpha Or Number Description||^[ \t]*(?<Index>[A-Z0-9])[\).:][ \t]+(?<Subject>[^:\r\n]+\r?\n(?:^[^ \r\n][^:\).][^:\r\n]+\r?\n)*)
