cancer link|tumor type|*body location|body location laterality|Pre-Diagnostic Start Date|Pre-Diagnostic End Date|Pre-Diagnostic Documents|Diagnostic Start Date|Diagnostic End Date|Diagnostic Documents|Treatment Start Date|Treatment End Date|Treatment Documents|Follow-up Start Date|Follow-up End Date|Follow-up Documentscancer_patientx_Left_Breast_Current|PrimaryTumor|Breast|Left|1/21/10|1/21/10|patientX_doc1_RAD.txt|1/30/10|1/30/10|patientX_doc2_SP.txt|12/2/10|12/2/10|patientX_doc3_NOTE.txt|||cancer_patientx_Left_Breast_Current|Regional_Metastasis|Axillary_Lymph_Node|Left|1/21/10|1/21/10|patientX_doc1_RAD.txt|1/30/10|1/30/10|patientX_doc2_SP.txt|12/2/10|12/2/10|patientX_doc3_NOTE.txt|||