-cancer ID|*patient ID|*body location|body location laterality|Temporality|clinical stage|clinical T classification|clinical N classification|clinical M classification|pathologic T classification|pathologic N classification|pathologic M classification|
cancer_patientX_Left_Breast_Current|patientX|Breast|Left|Current|Stage_2A|||||||
